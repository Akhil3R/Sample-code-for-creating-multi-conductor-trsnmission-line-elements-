* 10-wire PI Transmission Line Subcircuit Model

.SUBCKT TRANSMISSION_LINE in1 out1 in2 out2 in3 out3 in4 out4 in5 out5 in6 out6 in7 out7 in8 out8 in9 out9 in10 out10
R0_1 node0_0 node0_0_mid 6.559697e-02
L0_1 node0_0_mid node1_0 1.324593e-01
R0_2 node0_1 node0_1_mid 6.559697e-02
L0_2 node0_1_mid node1_1 1.324593e-01
R0_3 node0_2 node0_2_mid 6.559697e-02
L0_3 node0_2_mid node1_2 1.324592e-01
R0_4 node0_3 node0_3_mid 6.559697e-02
L0_4 node0_3_mid node1_3 1.324592e-01
R0_5 node0_4 node0_4_mid 6.559697e-02
L0_5 node0_4_mid node1_4 1.324592e-01
R0_6 node0_5 node0_5_mid 6.559697e-02
L0_6 node0_5_mid node1_5 1.324591e-01
R0_7 node0_6 node0_6_mid 6.559697e-02
L0_7 node0_6_mid node1_6 1.324591e-01
R0_8 node0_7 node0_7_mid 6.559697e-02
L0_8 node0_7_mid node1_7 1.324591e-01
R0_9 node0_8 node0_8_mid 6.559697e-02
L0_9 node0_8_mid node1_8 1.324591e-01
R0_10 node0_9 node0_9_mid 6.559697e-02
L0_10 node0_9_mid node1_9 1.324591e-01
K0_1 L0_1 L0_2 1.000000e+00
K0_2 L0_1 L0_3 1.000000e+00
K0_3 L0_1 L0_4 1.000000e+00
K0_4 L0_1 L0_5 1.000000e+00
K0_5 L0_1 L0_6 9.999999e-01
K0_6 L0_1 L0_7 1.000000e+00
K0_7 L0_1 L0_8 9.999999e-01
K0_8 L0_1 L0_9 9.999999e-01
K0_9 L0_1 L0_10 9.999999e-01
K0_10 L0_2 L0_3 1.000000e+00
K0_11 L0_2 L0_4 1.000000e+00
K0_12 L0_2 L0_5 1.000000e+00
K0_13 L0_2 L0_6 9.999999e-01
K0_14 L0_2 L0_7 1.000000e+00
K0_15 L0_2 L0_8 9.999999e-01
K0_16 L0_2 L0_9 9.999999e-01
K0_17 L0_2 L0_10 9.999999e-01
K0_18 L0_3 L0_4 1.000000e+00
K0_19 L0_3 L0_5 1.000000e+00
K0_20 L0_3 L0_6 9.999999e-01
K0_21 L0_3 L0_7 9.999999e-01
K0_22 L0_3 L0_8 9.999999e-01
K0_23 L0_3 L0_9 9.999999e-01
K0_24 L0_3 L0_10 9.999998e-01
K0_25 L0_4 L0_5 1.000000e+00
K0_26 L0_4 L0_6 9.999999e-01
K0_27 L0_4 L0_7 1.000000e+00
K0_28 L0_4 L0_8 9.999999e-01
K0_29 L0_4 L0_9 9.999999e-01
K0_30 L0_4 L0_10 9.999999e-01
K0_31 L0_5 L0_6 9.999999e-01
K0_32 L0_5 L0_7 1.000000e+00
K0_33 L0_5 L0_8 9.999999e-01
K0_34 L0_5 L0_9 9.999999e-01
K0_35 L0_5 L0_10 9.999999e-01
K0_36 L0_6 L0_7 9.999999e-01
K0_37 L0_6 L0_8 1.000000e+00
K0_38 L0_6 L0_9 1.000000e+00
K0_39 L0_6 L0_10 9.999999e-01
K0_40 L0_7 L0_8 9.999999e-01
K0_41 L0_7 L0_9 9.999999e-01
K0_42 L0_7 L0_10 9.999999e-01
K0_43 L0_8 L0_9 1.000000e+00
K0_44 L0_8 L0_10 1.000000e+00
K0_45 L0_9 L0_10 1.000000e+00
C0_1 node1_0 0 4.303416e-13
G0_1 node1_0 0 node1_0 0 2.703916e-06
C0_2 node1_1 0 6.975560e-13
G0_2 node1_1 0 node1_1 0 4.382874e-06
C0_3 node1_2 0 7.023171e-13
G0_3 node1_2 0 node1_2 0 4.412789e-06
C0_4 node1_3 0 7.031524e-13
G0_4 node1_3 0 node1_3 0 4.418037e-06
C0_5 node1_4 0 7.034466e-13
G0_5 node1_4 0 node1_4 0 4.419885e-06
C0_6 node1_5 0 7.035676e-13
G0_6 node1_5 0 node1_5 0 4.420645e-06
C0_7 node1_6 0 7.030741e-13
G0_7 node1_6 0 node1_6 0 4.417545e-06
C0_8 node1_7 0 7.018853e-13
G0_8 node1_7 0 node1_7 0 4.410075e-06
C0_9 node1_8 0 6.973380e-13
G0_9 node1_8 0 node1_8 0 4.381504e-06
C0_10 node1_9 0 4.303249e-13
G0_10 node1_9 0 node1_9 0 2.703811e-06
CM0_1 node1_0 node1_1 -3.372270e-13
CM0_2 node1_0 node1_2 -4.333637e-14
CM0_3 node1_0 node1_3 -2.097687e-14
CM0_4 node1_0 node1_4 -1.177420e-14
CM0_5 node1_0 node1_5 -6.918544e-15
CM0_6 node1_0 node1_6 -4.146150e-15
CM0_7 node1_0 node1_7 -2.537949e-15
CM0_8 node1_0 node1_8 -1.643541e-15
CM0_9 node1_0 node1_9 -1.780983e-15
CM0_10 node1_1 node1_2 -3.044883e-13
CM0_11 node1_1 node1_3 -2.759806e-14
CM0_12 node1_1 node1_4 -1.220281e-14
CM0_13 node1_1 node1_5 -6.645893e-15
CM0_14 node1_1 node1_6 -3.879486e-15
CM0_15 node1_1 node1_7 -2.352696e-15
CM0_16 node1_1 node1_8 -1.518489e-15
CM0_17 node1_1 node1_9 -1.643380e-15
CM0_18 node1_2 node1_3 -3.019823e-13
CM0_19 node1_2 node1_4 -2.628447e-14
CM0_20 node1_2 node1_5 -1.143815e-14
CM0_21 node1_2 node1_6 -6.217217e-15
CM0_22 node1_2 node1_7 -3.678469e-15
CM0_23 node1_2 node1_8 -2.353400e-15
CM0_24 node1_2 node1_9 -2.538483e-15
CM0_25 node1_3 node1_4 -3.011554e-13
CM0_26 node1_3 node1_5 -2.592703e-14
CM0_27 node1_3 node1_6 -1.127554e-14
CM0_28 node1_3 node1_7 -6.213871e-15
CM0_29 node1_3 node1_8 -3.878491e-15
CM0_30 node1_3 node1_9 -4.144789e-15
CM0_31 node1_4 node1_5 -3.011387e-13
CM0_32 node1_4 node1_6 -2.590566e-14
CM0_33 node1_4 node1_7 -1.142857e-14
CM0_34 node1_4 node1_8 -6.642276e-15
CM0_35 node1_4 node1_9 -6.914501e-15
CM0_36 node1_5 node1_6 -3.012291e-13
CM0_37 node1_5 node1_7 -2.628136e-14
CM0_38 node1_5 node1_8 -1.220907e-14
CM0_39 node1_5 node1_9 -1.177964e-14
CM0_40 node1_6 node1_7 -3.018016e-13
CM0_41 node1_6 node1_8 -2.762580e-14
CM0_42 node1_6 node1_9 -2.099353e-14
CM0_43 node1_7 node1_8 -3.042640e-13
CM0_44 node1_7 node1_9 -4.332676e-14
CM0_45 node1_8 node1_9 -3.372029e-13
R1_1 node1_0 node1_0_mid 6.559697e-02
L1_1 node1_0_mid node2_0 1.324593e-01
R1_2 node1_1 node1_1_mid 6.559697e-02
L1_2 node1_1_mid node2_1 1.324593e-01
R1_3 node1_2 node1_2_mid 6.559697e-02
L1_3 node1_2_mid node2_2 1.324592e-01
R1_4 node1_3 node1_3_mid 6.559697e-02
L1_4 node1_3_mid node2_3 1.324592e-01
R1_5 node1_4 node1_4_mid 6.559697e-02
L1_5 node1_4_mid node2_4 1.324592e-01
R1_6 node1_5 node1_5_mid 6.559697e-02
L1_6 node1_5_mid node2_5 1.324591e-01
R1_7 node1_6 node1_6_mid 6.559697e-02
L1_7 node1_6_mid node2_6 1.324591e-01
R1_8 node1_7 node1_7_mid 6.559697e-02
L1_8 node1_7_mid node2_7 1.324591e-01
R1_9 node1_8 node1_8_mid 6.559697e-02
L1_9 node1_8_mid node2_8 1.324591e-01
R1_10 node1_9 node1_9_mid 6.559697e-02
L1_10 node1_9_mid node2_9 1.324591e-01
K1_1 L1_1 L1_2 1.000000e+00
K1_2 L1_1 L1_3 1.000000e+00
K1_3 L1_1 L1_4 1.000000e+00
K1_4 L1_1 L1_5 1.000000e+00
K1_5 L1_1 L1_6 9.999999e-01
K1_6 L1_1 L1_7 1.000000e+00
K1_7 L1_1 L1_8 9.999999e-01
K1_8 L1_1 L1_9 9.999999e-01
K1_9 L1_1 L1_10 9.999999e-01
K1_10 L1_2 L1_3 1.000000e+00
K1_11 L1_2 L1_4 1.000000e+00
K1_12 L1_2 L1_5 1.000000e+00
K1_13 L1_2 L1_6 9.999999e-01
K1_14 L1_2 L1_7 1.000000e+00
K1_15 L1_2 L1_8 9.999999e-01
K1_16 L1_2 L1_9 9.999999e-01
K1_17 L1_2 L1_10 9.999999e-01
K1_18 L1_3 L1_4 1.000000e+00
K1_19 L1_3 L1_5 1.000000e+00
K1_20 L1_3 L1_6 9.999999e-01
K1_21 L1_3 L1_7 9.999999e-01
K1_22 L1_3 L1_8 9.999999e-01
K1_23 L1_3 L1_9 9.999999e-01
K1_24 L1_3 L1_10 9.999998e-01
K1_25 L1_4 L1_5 1.000000e+00
K1_26 L1_4 L1_6 9.999999e-01
K1_27 L1_4 L1_7 1.000000e+00
K1_28 L1_4 L1_8 9.999999e-01
K1_29 L1_4 L1_9 9.999999e-01
K1_30 L1_4 L1_10 9.999999e-01
K1_31 L1_5 L1_6 9.999999e-01
K1_32 L1_5 L1_7 1.000000e+00
K1_33 L1_5 L1_8 9.999999e-01
K1_34 L1_5 L1_9 9.999999e-01
K1_35 L1_5 L1_10 9.999999e-01
K1_36 L1_6 L1_7 9.999999e-01
K1_37 L1_6 L1_8 1.000000e+00
K1_38 L1_6 L1_9 1.000000e+00
K1_39 L1_6 L1_10 9.999999e-01
K1_40 L1_7 L1_8 9.999999e-01
K1_41 L1_7 L1_9 9.999999e-01
K1_42 L1_7 L1_10 9.999999e-01
K1_43 L1_8 L1_9 1.000000e+00
K1_44 L1_8 L1_10 1.000000e+00
K1_45 L1_9 L1_10 1.000000e+00
C1_1 node2_0 0 4.303416e-13
G1_1 node2_0 0 node2_0 0 2.703916e-06
C1_2 node2_1 0 6.975560e-13
G1_2 node2_1 0 node2_1 0 4.382874e-06
C1_3 node2_2 0 7.023171e-13
G1_3 node2_2 0 node2_2 0 4.412789e-06
C1_4 node2_3 0 7.031524e-13
G1_4 node2_3 0 node2_3 0 4.418037e-06
C1_5 node2_4 0 7.034466e-13
G1_5 node2_4 0 node2_4 0 4.419885e-06
C1_6 node2_5 0 7.035676e-13
G1_6 node2_5 0 node2_5 0 4.420645e-06
C1_7 node2_6 0 7.030741e-13
G1_7 node2_6 0 node2_6 0 4.417545e-06
C1_8 node2_7 0 7.018853e-13
G1_8 node2_7 0 node2_7 0 4.410075e-06
C1_9 node2_8 0 6.973380e-13
G1_9 node2_8 0 node2_8 0 4.381504e-06
C1_10 node2_9 0 4.303249e-13
G1_10 node2_9 0 node2_9 0 2.703811e-06
CM1_1 node2_0 node2_1 -3.372270e-13
CM1_2 node2_0 node2_2 -4.333637e-14
CM1_3 node2_0 node2_3 -2.097687e-14
CM1_4 node2_0 node2_4 -1.177420e-14
CM1_5 node2_0 node2_5 -6.918544e-15
CM1_6 node2_0 node2_6 -4.146150e-15
CM1_7 node2_0 node2_7 -2.537949e-15
CM1_8 node2_0 node2_8 -1.643541e-15
CM1_9 node2_0 node2_9 -1.780983e-15
CM1_10 node2_1 node2_2 -3.044883e-13
CM1_11 node2_1 node2_3 -2.759806e-14
CM1_12 node2_1 node2_4 -1.220281e-14
CM1_13 node2_1 node2_5 -6.645893e-15
CM1_14 node2_1 node2_6 -3.879486e-15
CM1_15 node2_1 node2_7 -2.352696e-15
CM1_16 node2_1 node2_8 -1.518489e-15
CM1_17 node2_1 node2_9 -1.643380e-15
CM1_18 node2_2 node2_3 -3.019823e-13
CM1_19 node2_2 node2_4 -2.628447e-14
CM1_20 node2_2 node2_5 -1.143815e-14
CM1_21 node2_2 node2_6 -6.217217e-15
CM1_22 node2_2 node2_7 -3.678469e-15
CM1_23 node2_2 node2_8 -2.353400e-15
CM1_24 node2_2 node2_9 -2.538483e-15
CM1_25 node2_3 node2_4 -3.011554e-13
CM1_26 node2_3 node2_5 -2.592703e-14
CM1_27 node2_3 node2_6 -1.127554e-14
CM1_28 node2_3 node2_7 -6.213871e-15
CM1_29 node2_3 node2_8 -3.878491e-15
CM1_30 node2_3 node2_9 -4.144789e-15
CM1_31 node2_4 node2_5 -3.011387e-13
CM1_32 node2_4 node2_6 -2.590566e-14
CM1_33 node2_4 node2_7 -1.142857e-14
CM1_34 node2_4 node2_8 -6.642276e-15
CM1_35 node2_4 node2_9 -6.914501e-15
CM1_36 node2_5 node2_6 -3.012291e-13
CM1_37 node2_5 node2_7 -2.628136e-14
CM1_38 node2_5 node2_8 -1.220907e-14
CM1_39 node2_5 node2_9 -1.177964e-14
CM1_40 node2_6 node2_7 -3.018016e-13
CM1_41 node2_6 node2_8 -2.762580e-14
CM1_42 node2_6 node2_9 -2.099353e-14
CM1_43 node2_7 node2_8 -3.042640e-13
CM1_44 node2_7 node2_9 -4.332676e-14
CM1_45 node2_8 node2_9 -3.372029e-13
R2_1 node2_0 node2_0_mid 6.559697e-02
L2_1 node2_0_mid node3_0 1.324593e-01
R2_2 node2_1 node2_1_mid 6.559697e-02
L2_2 node2_1_mid node3_1 1.324593e-01
R2_3 node2_2 node2_2_mid 6.559697e-02
L2_3 node2_2_mid node3_2 1.324592e-01
R2_4 node2_3 node2_3_mid 6.559697e-02
L2_4 node2_3_mid node3_3 1.324592e-01
R2_5 node2_4 node2_4_mid 6.559697e-02
L2_5 node2_4_mid node3_4 1.324592e-01
R2_6 node2_5 node2_5_mid 6.559697e-02
L2_6 node2_5_mid node3_5 1.324591e-01
R2_7 node2_6 node2_6_mid 6.559697e-02
L2_7 node2_6_mid node3_6 1.324591e-01
R2_8 node2_7 node2_7_mid 6.559697e-02
L2_8 node2_7_mid node3_7 1.324591e-01
R2_9 node2_8 node2_8_mid 6.559697e-02
L2_9 node2_8_mid node3_8 1.324591e-01
R2_10 node2_9 node2_9_mid 6.559697e-02
L2_10 node2_9_mid node3_9 1.324591e-01
K2_1 L2_1 L2_2 1.000000e+00
K2_2 L2_1 L2_3 1.000000e+00
K2_3 L2_1 L2_4 1.000000e+00
K2_4 L2_1 L2_5 1.000000e+00
K2_5 L2_1 L2_6 9.999999e-01
K2_6 L2_1 L2_7 1.000000e+00
K2_7 L2_1 L2_8 9.999999e-01
K2_8 L2_1 L2_9 9.999999e-01
K2_9 L2_1 L2_10 9.999999e-01
K2_10 L2_2 L2_3 1.000000e+00
K2_11 L2_2 L2_4 1.000000e+00
K2_12 L2_2 L2_5 1.000000e+00
K2_13 L2_2 L2_6 9.999999e-01
K2_14 L2_2 L2_7 1.000000e+00
K2_15 L2_2 L2_8 9.999999e-01
K2_16 L2_2 L2_9 9.999999e-01
K2_17 L2_2 L2_10 9.999999e-01
K2_18 L2_3 L2_4 1.000000e+00
K2_19 L2_3 L2_5 1.000000e+00
K2_20 L2_3 L2_6 9.999999e-01
K2_21 L2_3 L2_7 9.999999e-01
K2_22 L2_3 L2_8 9.999999e-01
K2_23 L2_3 L2_9 9.999999e-01
K2_24 L2_3 L2_10 9.999998e-01
K2_25 L2_4 L2_5 1.000000e+00
K2_26 L2_4 L2_6 9.999999e-01
K2_27 L2_4 L2_7 1.000000e+00
K2_28 L2_4 L2_8 9.999999e-01
K2_29 L2_4 L2_9 9.999999e-01
K2_30 L2_4 L2_10 9.999999e-01
K2_31 L2_5 L2_6 9.999999e-01
K2_32 L2_5 L2_7 1.000000e+00
K2_33 L2_5 L2_8 9.999999e-01
K2_34 L2_5 L2_9 9.999999e-01
K2_35 L2_5 L2_10 9.999999e-01
K2_36 L2_6 L2_7 9.999999e-01
K2_37 L2_6 L2_8 1.000000e+00
K2_38 L2_6 L2_9 1.000000e+00
K2_39 L2_6 L2_10 9.999999e-01
K2_40 L2_7 L2_8 9.999999e-01
K2_41 L2_7 L2_9 9.999999e-01
K2_42 L2_7 L2_10 9.999999e-01
K2_43 L2_8 L2_9 1.000000e+00
K2_44 L2_8 L2_10 1.000000e+00
K2_45 L2_9 L2_10 1.000000e+00
C2_1 node3_0 0 4.303416e-13
G2_1 node3_0 0 node3_0 0 2.703916e-06
C2_2 node3_1 0 6.975560e-13
G2_2 node3_1 0 node3_1 0 4.382874e-06
C2_3 node3_2 0 7.023171e-13
G2_3 node3_2 0 node3_2 0 4.412789e-06
C2_4 node3_3 0 7.031524e-13
G2_4 node3_3 0 node3_3 0 4.418037e-06
C2_5 node3_4 0 7.034466e-13
G2_5 node3_4 0 node3_4 0 4.419885e-06
C2_6 node3_5 0 7.035676e-13
G2_6 node3_5 0 node3_5 0 4.420645e-06
C2_7 node3_6 0 7.030741e-13
G2_7 node3_6 0 node3_6 0 4.417545e-06
C2_8 node3_7 0 7.018853e-13
G2_8 node3_7 0 node3_7 0 4.410075e-06
C2_9 node3_8 0 6.973380e-13
G2_9 node3_8 0 node3_8 0 4.381504e-06
C2_10 node3_9 0 4.303249e-13
G2_10 node3_9 0 node3_9 0 2.703811e-06
CM2_1 node3_0 node3_1 -3.372270e-13
CM2_2 node3_0 node3_2 -4.333637e-14
CM2_3 node3_0 node3_3 -2.097687e-14
CM2_4 node3_0 node3_4 -1.177420e-14
CM2_5 node3_0 node3_5 -6.918544e-15
CM2_6 node3_0 node3_6 -4.146150e-15
CM2_7 node3_0 node3_7 -2.537949e-15
CM2_8 node3_0 node3_8 -1.643541e-15
CM2_9 node3_0 node3_9 -1.780983e-15
CM2_10 node3_1 node3_2 -3.044883e-13
CM2_11 node3_1 node3_3 -2.759806e-14
CM2_12 node3_1 node3_4 -1.220281e-14
CM2_13 node3_1 node3_5 -6.645893e-15
CM2_14 node3_1 node3_6 -3.879486e-15
CM2_15 node3_1 node3_7 -2.352696e-15
CM2_16 node3_1 node3_8 -1.518489e-15
CM2_17 node3_1 node3_9 -1.643380e-15
CM2_18 node3_2 node3_3 -3.019823e-13
CM2_19 node3_2 node3_4 -2.628447e-14
CM2_20 node3_2 node3_5 -1.143815e-14
CM2_21 node3_2 node3_6 -6.217217e-15
CM2_22 node3_2 node3_7 -3.678469e-15
CM2_23 node3_2 node3_8 -2.353400e-15
CM2_24 node3_2 node3_9 -2.538483e-15
CM2_25 node3_3 node3_4 -3.011554e-13
CM2_26 node3_3 node3_5 -2.592703e-14
CM2_27 node3_3 node3_6 -1.127554e-14
CM2_28 node3_3 node3_7 -6.213871e-15
CM2_29 node3_3 node3_8 -3.878491e-15
CM2_30 node3_3 node3_9 -4.144789e-15
CM2_31 node3_4 node3_5 -3.011387e-13
CM2_32 node3_4 node3_6 -2.590566e-14
CM2_33 node3_4 node3_7 -1.142857e-14
CM2_34 node3_4 node3_8 -6.642276e-15
CM2_35 node3_4 node3_9 -6.914501e-15
CM2_36 node3_5 node3_6 -3.012291e-13
CM2_37 node3_5 node3_7 -2.628136e-14
CM2_38 node3_5 node3_8 -1.220907e-14
CM2_39 node3_5 node3_9 -1.177964e-14
CM2_40 node3_6 node3_7 -3.018016e-13
CM2_41 node3_6 node3_8 -2.762580e-14
CM2_42 node3_6 node3_9 -2.099353e-14
CM2_43 node3_7 node3_8 -3.042640e-13
CM2_44 node3_7 node3_9 -4.332676e-14
CM2_45 node3_8 node3_9 -3.372029e-13
R3_1 node3_0 node3_0_mid 6.559697e-02
L3_1 node3_0_mid node4_0 1.324593e-01
R3_2 node3_1 node3_1_mid 6.559697e-02
L3_2 node3_1_mid node4_1 1.324593e-01
R3_3 node3_2 node3_2_mid 6.559697e-02
L3_3 node3_2_mid node4_2 1.324592e-01
R3_4 node3_3 node3_3_mid 6.559697e-02
L3_4 node3_3_mid node4_3 1.324592e-01
R3_5 node3_4 node3_4_mid 6.559697e-02
L3_5 node3_4_mid node4_4 1.324592e-01
R3_6 node3_5 node3_5_mid 6.559697e-02
L3_6 node3_5_mid node4_5 1.324591e-01
R3_7 node3_6 node3_6_mid 6.559697e-02
L3_7 node3_6_mid node4_6 1.324591e-01
R3_8 node3_7 node3_7_mid 6.559697e-02
L3_8 node3_7_mid node4_7 1.324591e-01
R3_9 node3_8 node3_8_mid 6.559697e-02
L3_9 node3_8_mid node4_8 1.324591e-01
R3_10 node3_9 node3_9_mid 6.559697e-02
L3_10 node3_9_mid node4_9 1.324591e-01
K3_1 L3_1 L3_2 1.000000e+00
K3_2 L3_1 L3_3 1.000000e+00
K3_3 L3_1 L3_4 1.000000e+00
K3_4 L3_1 L3_5 1.000000e+00
K3_5 L3_1 L3_6 9.999999e-01
K3_6 L3_1 L3_7 1.000000e+00
K3_7 L3_1 L3_8 9.999999e-01
K3_8 L3_1 L3_9 9.999999e-01
K3_9 L3_1 L3_10 9.999999e-01
K3_10 L3_2 L3_3 1.000000e+00
K3_11 L3_2 L3_4 1.000000e+00
K3_12 L3_2 L3_5 1.000000e+00
K3_13 L3_2 L3_6 9.999999e-01
K3_14 L3_2 L3_7 1.000000e+00
K3_15 L3_2 L3_8 9.999999e-01
K3_16 L3_2 L3_9 9.999999e-01
K3_17 L3_2 L3_10 9.999999e-01
K3_18 L3_3 L3_4 1.000000e+00
K3_19 L3_3 L3_5 1.000000e+00
K3_20 L3_3 L3_6 9.999999e-01
K3_21 L3_3 L3_7 9.999999e-01
K3_22 L3_3 L3_8 9.999999e-01
K3_23 L3_3 L3_9 9.999999e-01
K3_24 L3_3 L3_10 9.999998e-01
K3_25 L3_4 L3_5 1.000000e+00
K3_26 L3_4 L3_6 9.999999e-01
K3_27 L3_4 L3_7 1.000000e+00
K3_28 L3_4 L3_8 9.999999e-01
K3_29 L3_4 L3_9 9.999999e-01
K3_30 L3_4 L3_10 9.999999e-01
K3_31 L3_5 L3_6 9.999999e-01
K3_32 L3_5 L3_7 1.000000e+00
K3_33 L3_5 L3_8 9.999999e-01
K3_34 L3_5 L3_9 9.999999e-01
K3_35 L3_5 L3_10 9.999999e-01
K3_36 L3_6 L3_7 9.999999e-01
K3_37 L3_6 L3_8 1.000000e+00
K3_38 L3_6 L3_9 1.000000e+00
K3_39 L3_6 L3_10 9.999999e-01
K3_40 L3_7 L3_8 9.999999e-01
K3_41 L3_7 L3_9 9.999999e-01
K3_42 L3_7 L3_10 9.999999e-01
K3_43 L3_8 L3_9 1.000000e+00
K3_44 L3_8 L3_10 1.000000e+00
K3_45 L3_9 L3_10 1.000000e+00
C3_1 node4_0 0 4.303416e-13
G3_1 node4_0 0 node4_0 0 2.703916e-06
C3_2 node4_1 0 6.975560e-13
G3_2 node4_1 0 node4_1 0 4.382874e-06
C3_3 node4_2 0 7.023171e-13
G3_3 node4_2 0 node4_2 0 4.412789e-06
C3_4 node4_3 0 7.031524e-13
G3_4 node4_3 0 node4_3 0 4.418037e-06
C3_5 node4_4 0 7.034466e-13
G3_5 node4_4 0 node4_4 0 4.419885e-06
C3_6 node4_5 0 7.035676e-13
G3_6 node4_5 0 node4_5 0 4.420645e-06
C3_7 node4_6 0 7.030741e-13
G3_7 node4_6 0 node4_6 0 4.417545e-06
C3_8 node4_7 0 7.018853e-13
G3_8 node4_7 0 node4_7 0 4.410075e-06
C3_9 node4_8 0 6.973380e-13
G3_9 node4_8 0 node4_8 0 4.381504e-06
C3_10 node4_9 0 4.303249e-13
G3_10 node4_9 0 node4_9 0 2.703811e-06
CM3_1 node4_0 node4_1 -3.372270e-13
CM3_2 node4_0 node4_2 -4.333637e-14
CM3_3 node4_0 node4_3 -2.097687e-14
CM3_4 node4_0 node4_4 -1.177420e-14
CM3_5 node4_0 node4_5 -6.918544e-15
CM3_6 node4_0 node4_6 -4.146150e-15
CM3_7 node4_0 node4_7 -2.537949e-15
CM3_8 node4_0 node4_8 -1.643541e-15
CM3_9 node4_0 node4_9 -1.780983e-15
CM3_10 node4_1 node4_2 -3.044883e-13
CM3_11 node4_1 node4_3 -2.759806e-14
CM3_12 node4_1 node4_4 -1.220281e-14
CM3_13 node4_1 node4_5 -6.645893e-15
CM3_14 node4_1 node4_6 -3.879486e-15
CM3_15 node4_1 node4_7 -2.352696e-15
CM3_16 node4_1 node4_8 -1.518489e-15
CM3_17 node4_1 node4_9 -1.643380e-15
CM3_18 node4_2 node4_3 -3.019823e-13
CM3_19 node4_2 node4_4 -2.628447e-14
CM3_20 node4_2 node4_5 -1.143815e-14
CM3_21 node4_2 node4_6 -6.217217e-15
CM3_22 node4_2 node4_7 -3.678469e-15
CM3_23 node4_2 node4_8 -2.353400e-15
CM3_24 node4_2 node4_9 -2.538483e-15
CM3_25 node4_3 node4_4 -3.011554e-13
CM3_26 node4_3 node4_5 -2.592703e-14
CM3_27 node4_3 node4_6 -1.127554e-14
CM3_28 node4_3 node4_7 -6.213871e-15
CM3_29 node4_3 node4_8 -3.878491e-15
CM3_30 node4_3 node4_9 -4.144789e-15
CM3_31 node4_4 node4_5 -3.011387e-13
CM3_32 node4_4 node4_6 -2.590566e-14
CM3_33 node4_4 node4_7 -1.142857e-14
CM3_34 node4_4 node4_8 -6.642276e-15
CM3_35 node4_4 node4_9 -6.914501e-15
CM3_36 node4_5 node4_6 -3.012291e-13
CM3_37 node4_5 node4_7 -2.628136e-14
CM3_38 node4_5 node4_8 -1.220907e-14
CM3_39 node4_5 node4_9 -1.177964e-14
CM3_40 node4_6 node4_7 -3.018016e-13
CM3_41 node4_6 node4_8 -2.762580e-14
CM3_42 node4_6 node4_9 -2.099353e-14
CM3_43 node4_7 node4_8 -3.042640e-13
CM3_44 node4_7 node4_9 -4.332676e-14
CM3_45 node4_8 node4_9 -3.372029e-13
R4_1 node4_0 node4_0_mid 6.559697e-02
L4_1 node4_0_mid node5_0 1.324593e-01
R4_2 node4_1 node4_1_mid 6.559697e-02
L4_2 node4_1_mid node5_1 1.324593e-01
R4_3 node4_2 node4_2_mid 6.559697e-02
L4_3 node4_2_mid node5_2 1.324592e-01
R4_4 node4_3 node4_3_mid 6.559697e-02
L4_4 node4_3_mid node5_3 1.324592e-01
R4_5 node4_4 node4_4_mid 6.559697e-02
L4_5 node4_4_mid node5_4 1.324592e-01
R4_6 node4_5 node4_5_mid 6.559697e-02
L4_6 node4_5_mid node5_5 1.324591e-01
R4_7 node4_6 node4_6_mid 6.559697e-02
L4_7 node4_6_mid node5_6 1.324591e-01
R4_8 node4_7 node4_7_mid 6.559697e-02
L4_8 node4_7_mid node5_7 1.324591e-01
R4_9 node4_8 node4_8_mid 6.559697e-02
L4_9 node4_8_mid node5_8 1.324591e-01
R4_10 node4_9 node4_9_mid 6.559697e-02
L4_10 node4_9_mid node5_9 1.324591e-01
K4_1 L4_1 L4_2 1.000000e+00
K4_2 L4_1 L4_3 1.000000e+00
K4_3 L4_1 L4_4 1.000000e+00
K4_4 L4_1 L4_5 1.000000e+00
K4_5 L4_1 L4_6 9.999999e-01
K4_6 L4_1 L4_7 1.000000e+00
K4_7 L4_1 L4_8 9.999999e-01
K4_8 L4_1 L4_9 9.999999e-01
K4_9 L4_1 L4_10 9.999999e-01
K4_10 L4_2 L4_3 1.000000e+00
K4_11 L4_2 L4_4 1.000000e+00
K4_12 L4_2 L4_5 1.000000e+00
K4_13 L4_2 L4_6 9.999999e-01
K4_14 L4_2 L4_7 1.000000e+00
K4_15 L4_2 L4_8 9.999999e-01
K4_16 L4_2 L4_9 9.999999e-01
K4_17 L4_2 L4_10 9.999999e-01
K4_18 L4_3 L4_4 1.000000e+00
K4_19 L4_3 L4_5 1.000000e+00
K4_20 L4_3 L4_6 9.999999e-01
K4_21 L4_3 L4_7 9.999999e-01
K4_22 L4_3 L4_8 9.999999e-01
K4_23 L4_3 L4_9 9.999999e-01
K4_24 L4_3 L4_10 9.999998e-01
K4_25 L4_4 L4_5 1.000000e+00
K4_26 L4_4 L4_6 9.999999e-01
K4_27 L4_4 L4_7 1.000000e+00
K4_28 L4_4 L4_8 9.999999e-01
K4_29 L4_4 L4_9 9.999999e-01
K4_30 L4_4 L4_10 9.999999e-01
K4_31 L4_5 L4_6 9.999999e-01
K4_32 L4_5 L4_7 1.000000e+00
K4_33 L4_5 L4_8 9.999999e-01
K4_34 L4_5 L4_9 9.999999e-01
K4_35 L4_5 L4_10 9.999999e-01
K4_36 L4_6 L4_7 9.999999e-01
K4_37 L4_6 L4_8 1.000000e+00
K4_38 L4_6 L4_9 1.000000e+00
K4_39 L4_6 L4_10 9.999999e-01
K4_40 L4_7 L4_8 9.999999e-01
K4_41 L4_7 L4_9 9.999999e-01
K4_42 L4_7 L4_10 9.999999e-01
K4_43 L4_8 L4_9 1.000000e+00
K4_44 L4_8 L4_10 1.000000e+00
K4_45 L4_9 L4_10 1.000000e+00
C4_1 node5_0 0 4.303416e-13
G4_1 node5_0 0 node5_0 0 2.703916e-06
C4_2 node5_1 0 6.975560e-13
G4_2 node5_1 0 node5_1 0 4.382874e-06
C4_3 node5_2 0 7.023171e-13
G4_3 node5_2 0 node5_2 0 4.412789e-06
C4_4 node5_3 0 7.031524e-13
G4_4 node5_3 0 node5_3 0 4.418037e-06
C4_5 node5_4 0 7.034466e-13
G4_5 node5_4 0 node5_4 0 4.419885e-06
C4_6 node5_5 0 7.035676e-13
G4_6 node5_5 0 node5_5 0 4.420645e-06
C4_7 node5_6 0 7.030741e-13
G4_7 node5_6 0 node5_6 0 4.417545e-06
C4_8 node5_7 0 7.018853e-13
G4_8 node5_7 0 node5_7 0 4.410075e-06
C4_9 node5_8 0 6.973380e-13
G4_9 node5_8 0 node5_8 0 4.381504e-06
C4_10 node5_9 0 4.303249e-13
G4_10 node5_9 0 node5_9 0 2.703811e-06
CM4_1 node5_0 node5_1 -3.372270e-13
CM4_2 node5_0 node5_2 -4.333637e-14
CM4_3 node5_0 node5_3 -2.097687e-14
CM4_4 node5_0 node5_4 -1.177420e-14
CM4_5 node5_0 node5_5 -6.918544e-15
CM4_6 node5_0 node5_6 -4.146150e-15
CM4_7 node5_0 node5_7 -2.537949e-15
CM4_8 node5_0 node5_8 -1.643541e-15
CM4_9 node5_0 node5_9 -1.780983e-15
CM4_10 node5_1 node5_2 -3.044883e-13
CM4_11 node5_1 node5_3 -2.759806e-14
CM4_12 node5_1 node5_4 -1.220281e-14
CM4_13 node5_1 node5_5 -6.645893e-15
CM4_14 node5_1 node5_6 -3.879486e-15
CM4_15 node5_1 node5_7 -2.352696e-15
CM4_16 node5_1 node5_8 -1.518489e-15
CM4_17 node5_1 node5_9 -1.643380e-15
CM4_18 node5_2 node5_3 -3.019823e-13
CM4_19 node5_2 node5_4 -2.628447e-14
CM4_20 node5_2 node5_5 -1.143815e-14
CM4_21 node5_2 node5_6 -6.217217e-15
CM4_22 node5_2 node5_7 -3.678469e-15
CM4_23 node5_2 node5_8 -2.353400e-15
CM4_24 node5_2 node5_9 -2.538483e-15
CM4_25 node5_3 node5_4 -3.011554e-13
CM4_26 node5_3 node5_5 -2.592703e-14
CM4_27 node5_3 node5_6 -1.127554e-14
CM4_28 node5_3 node5_7 -6.213871e-15
CM4_29 node5_3 node5_8 -3.878491e-15
CM4_30 node5_3 node5_9 -4.144789e-15
CM4_31 node5_4 node5_5 -3.011387e-13
CM4_32 node5_4 node5_6 -2.590566e-14
CM4_33 node5_4 node5_7 -1.142857e-14
CM4_34 node5_4 node5_8 -6.642276e-15
CM4_35 node5_4 node5_9 -6.914501e-15
CM4_36 node5_5 node5_6 -3.012291e-13
CM4_37 node5_5 node5_7 -2.628136e-14
CM4_38 node5_5 node5_8 -1.220907e-14
CM4_39 node5_5 node5_9 -1.177964e-14
CM4_40 node5_6 node5_7 -3.018016e-13
CM4_41 node5_6 node5_8 -2.762580e-14
CM4_42 node5_6 node5_9 -2.099353e-14
CM4_43 node5_7 node5_8 -3.042640e-13
CM4_44 node5_7 node5_9 -4.332676e-14
CM4_45 node5_8 node5_9 -3.372029e-13
R5_1 node5_0 node5_0_mid 6.559697e-02
L5_1 node5_0_mid node6_0 1.324593e-01
R5_2 node5_1 node5_1_mid 6.559697e-02
L5_2 node5_1_mid node6_1 1.324593e-01
R5_3 node5_2 node5_2_mid 6.559697e-02
L5_3 node5_2_mid node6_2 1.324592e-01
R5_4 node5_3 node5_3_mid 6.559697e-02
L5_4 node5_3_mid node6_3 1.324592e-01
R5_5 node5_4 node5_4_mid 6.559697e-02
L5_5 node5_4_mid node6_4 1.324592e-01
R5_6 node5_5 node5_5_mid 6.559697e-02
L5_6 node5_5_mid node6_5 1.324591e-01
R5_7 node5_6 node5_6_mid 6.559697e-02
L5_7 node5_6_mid node6_6 1.324591e-01
R5_8 node5_7 node5_7_mid 6.559697e-02
L5_8 node5_7_mid node6_7 1.324591e-01
R5_9 node5_8 node5_8_mid 6.559697e-02
L5_9 node5_8_mid node6_8 1.324591e-01
R5_10 node5_9 node5_9_mid 6.559697e-02
L5_10 node5_9_mid node6_9 1.324591e-01
K5_1 L5_1 L5_2 1.000000e+00
K5_2 L5_1 L5_3 1.000000e+00
K5_3 L5_1 L5_4 1.000000e+00
K5_4 L5_1 L5_5 1.000000e+00
K5_5 L5_1 L5_6 9.999999e-01
K5_6 L5_1 L5_7 1.000000e+00
K5_7 L5_1 L5_8 9.999999e-01
K5_8 L5_1 L5_9 9.999999e-01
K5_9 L5_1 L5_10 9.999999e-01
K5_10 L5_2 L5_3 1.000000e+00
K5_11 L5_2 L5_4 1.000000e+00
K5_12 L5_2 L5_5 1.000000e+00
K5_13 L5_2 L5_6 9.999999e-01
K5_14 L5_2 L5_7 1.000000e+00
K5_15 L5_2 L5_8 9.999999e-01
K5_16 L5_2 L5_9 9.999999e-01
K5_17 L5_2 L5_10 9.999999e-01
K5_18 L5_3 L5_4 1.000000e+00
K5_19 L5_3 L5_5 1.000000e+00
K5_20 L5_3 L5_6 9.999999e-01
K5_21 L5_3 L5_7 9.999999e-01
K5_22 L5_3 L5_8 9.999999e-01
K5_23 L5_3 L5_9 9.999999e-01
K5_24 L5_3 L5_10 9.999998e-01
K5_25 L5_4 L5_5 1.000000e+00
K5_26 L5_4 L5_6 9.999999e-01
K5_27 L5_4 L5_7 1.000000e+00
K5_28 L5_4 L5_8 9.999999e-01
K5_29 L5_4 L5_9 9.999999e-01
K5_30 L5_4 L5_10 9.999999e-01
K5_31 L5_5 L5_6 9.999999e-01
K5_32 L5_5 L5_7 1.000000e+00
K5_33 L5_5 L5_8 9.999999e-01
K5_34 L5_5 L5_9 9.999999e-01
K5_35 L5_5 L5_10 9.999999e-01
K5_36 L5_6 L5_7 9.999999e-01
K5_37 L5_6 L5_8 1.000000e+00
K5_38 L5_6 L5_9 1.000000e+00
K5_39 L5_6 L5_10 9.999999e-01
K5_40 L5_7 L5_8 9.999999e-01
K5_41 L5_7 L5_9 9.999999e-01
K5_42 L5_7 L5_10 9.999999e-01
K5_43 L5_8 L5_9 1.000000e+00
K5_44 L5_8 L5_10 1.000000e+00
K5_45 L5_9 L5_10 1.000000e+00
C5_1 node6_0 0 4.303416e-13
G5_1 node6_0 0 node6_0 0 2.703916e-06
C5_2 node6_1 0 6.975560e-13
G5_2 node6_1 0 node6_1 0 4.382874e-06
C5_3 node6_2 0 7.023171e-13
G5_3 node6_2 0 node6_2 0 4.412789e-06
C5_4 node6_3 0 7.031524e-13
G5_4 node6_3 0 node6_3 0 4.418037e-06
C5_5 node6_4 0 7.034466e-13
G5_5 node6_4 0 node6_4 0 4.419885e-06
C5_6 node6_5 0 7.035676e-13
G5_6 node6_5 0 node6_5 0 4.420645e-06
C5_7 node6_6 0 7.030741e-13
G5_7 node6_6 0 node6_6 0 4.417545e-06
C5_8 node6_7 0 7.018853e-13
G5_8 node6_7 0 node6_7 0 4.410075e-06
C5_9 node6_8 0 6.973380e-13
G5_9 node6_8 0 node6_8 0 4.381504e-06
C5_10 node6_9 0 4.303249e-13
G5_10 node6_9 0 node6_9 0 2.703811e-06
CM5_1 node6_0 node6_1 -3.372270e-13
CM5_2 node6_0 node6_2 -4.333637e-14
CM5_3 node6_0 node6_3 -2.097687e-14
CM5_4 node6_0 node6_4 -1.177420e-14
CM5_5 node6_0 node6_5 -6.918544e-15
CM5_6 node6_0 node6_6 -4.146150e-15
CM5_7 node6_0 node6_7 -2.537949e-15
CM5_8 node6_0 node6_8 -1.643541e-15
CM5_9 node6_0 node6_9 -1.780983e-15
CM5_10 node6_1 node6_2 -3.044883e-13
CM5_11 node6_1 node6_3 -2.759806e-14
CM5_12 node6_1 node6_4 -1.220281e-14
CM5_13 node6_1 node6_5 -6.645893e-15
CM5_14 node6_1 node6_6 -3.879486e-15
CM5_15 node6_1 node6_7 -2.352696e-15
CM5_16 node6_1 node6_8 -1.518489e-15
CM5_17 node6_1 node6_9 -1.643380e-15
CM5_18 node6_2 node6_3 -3.019823e-13
CM5_19 node6_2 node6_4 -2.628447e-14
CM5_20 node6_2 node6_5 -1.143815e-14
CM5_21 node6_2 node6_6 -6.217217e-15
CM5_22 node6_2 node6_7 -3.678469e-15
CM5_23 node6_2 node6_8 -2.353400e-15
CM5_24 node6_2 node6_9 -2.538483e-15
CM5_25 node6_3 node6_4 -3.011554e-13
CM5_26 node6_3 node6_5 -2.592703e-14
CM5_27 node6_3 node6_6 -1.127554e-14
CM5_28 node6_3 node6_7 -6.213871e-15
CM5_29 node6_3 node6_8 -3.878491e-15
CM5_30 node6_3 node6_9 -4.144789e-15
CM5_31 node6_4 node6_5 -3.011387e-13
CM5_32 node6_4 node6_6 -2.590566e-14
CM5_33 node6_4 node6_7 -1.142857e-14
CM5_34 node6_4 node6_8 -6.642276e-15
CM5_35 node6_4 node6_9 -6.914501e-15
CM5_36 node6_5 node6_6 -3.012291e-13
CM5_37 node6_5 node6_7 -2.628136e-14
CM5_38 node6_5 node6_8 -1.220907e-14
CM5_39 node6_5 node6_9 -1.177964e-14
CM5_40 node6_6 node6_7 -3.018016e-13
CM5_41 node6_6 node6_8 -2.762580e-14
CM5_42 node6_6 node6_9 -2.099353e-14
CM5_43 node6_7 node6_8 -3.042640e-13
CM5_44 node6_7 node6_9 -4.332676e-14
CM5_45 node6_8 node6_9 -3.372029e-13
R6_1 node6_0 node6_0_mid 6.559697e-02
L6_1 node6_0_mid node7_0 1.324593e-01
R6_2 node6_1 node6_1_mid 6.559697e-02
L6_2 node6_1_mid node7_1 1.324593e-01
R6_3 node6_2 node6_2_mid 6.559697e-02
L6_3 node6_2_mid node7_2 1.324592e-01
R6_4 node6_3 node6_3_mid 6.559697e-02
L6_4 node6_3_mid node7_3 1.324592e-01
R6_5 node6_4 node6_4_mid 6.559697e-02
L6_5 node6_4_mid node7_4 1.324592e-01
R6_6 node6_5 node6_5_mid 6.559697e-02
L6_6 node6_5_mid node7_5 1.324591e-01
R6_7 node6_6 node6_6_mid 6.559697e-02
L6_7 node6_6_mid node7_6 1.324591e-01
R6_8 node6_7 node6_7_mid 6.559697e-02
L6_8 node6_7_mid node7_7 1.324591e-01
R6_9 node6_8 node6_8_mid 6.559697e-02
L6_9 node6_8_mid node7_8 1.324591e-01
R6_10 node6_9 node6_9_mid 6.559697e-02
L6_10 node6_9_mid node7_9 1.324591e-01
K6_1 L6_1 L6_2 1.000000e+00
K6_2 L6_1 L6_3 1.000000e+00
K6_3 L6_1 L6_4 1.000000e+00
K6_4 L6_1 L6_5 1.000000e+00
K6_5 L6_1 L6_6 9.999999e-01
K6_6 L6_1 L6_7 1.000000e+00
K6_7 L6_1 L6_8 9.999999e-01
K6_8 L6_1 L6_9 9.999999e-01
K6_9 L6_1 L6_10 9.999999e-01
K6_10 L6_2 L6_3 1.000000e+00
K6_11 L6_2 L6_4 1.000000e+00
K6_12 L6_2 L6_5 1.000000e+00
K6_13 L6_2 L6_6 9.999999e-01
K6_14 L6_2 L6_7 1.000000e+00
K6_15 L6_2 L6_8 9.999999e-01
K6_16 L6_2 L6_9 9.999999e-01
K6_17 L6_2 L6_10 9.999999e-01
K6_18 L6_3 L6_4 1.000000e+00
K6_19 L6_3 L6_5 1.000000e+00
K6_20 L6_3 L6_6 9.999999e-01
K6_21 L6_3 L6_7 9.999999e-01
K6_22 L6_3 L6_8 9.999999e-01
K6_23 L6_3 L6_9 9.999999e-01
K6_24 L6_3 L6_10 9.999998e-01
K6_25 L6_4 L6_5 1.000000e+00
K6_26 L6_4 L6_6 9.999999e-01
K6_27 L6_4 L6_7 1.000000e+00
K6_28 L6_4 L6_8 9.999999e-01
K6_29 L6_4 L6_9 9.999999e-01
K6_30 L6_4 L6_10 9.999999e-01
K6_31 L6_5 L6_6 9.999999e-01
K6_32 L6_5 L6_7 1.000000e+00
K6_33 L6_5 L6_8 9.999999e-01
K6_34 L6_5 L6_9 9.999999e-01
K6_35 L6_5 L6_10 9.999999e-01
K6_36 L6_6 L6_7 9.999999e-01
K6_37 L6_6 L6_8 1.000000e+00
K6_38 L6_6 L6_9 1.000000e+00
K6_39 L6_6 L6_10 9.999999e-01
K6_40 L6_7 L6_8 9.999999e-01
K6_41 L6_7 L6_9 9.999999e-01
K6_42 L6_7 L6_10 9.999999e-01
K6_43 L6_8 L6_9 1.000000e+00
K6_44 L6_8 L6_10 1.000000e+00
K6_45 L6_9 L6_10 1.000000e+00
C6_1 node7_0 0 4.303416e-13
G6_1 node7_0 0 node7_0 0 2.703916e-06
C6_2 node7_1 0 6.975560e-13
G6_2 node7_1 0 node7_1 0 4.382874e-06
C6_3 node7_2 0 7.023171e-13
G6_3 node7_2 0 node7_2 0 4.412789e-06
C6_4 node7_3 0 7.031524e-13
G6_4 node7_3 0 node7_3 0 4.418037e-06
C6_5 node7_4 0 7.034466e-13
G6_5 node7_4 0 node7_4 0 4.419885e-06
C6_6 node7_5 0 7.035676e-13
G6_6 node7_5 0 node7_5 0 4.420645e-06
C6_7 node7_6 0 7.030741e-13
G6_7 node7_6 0 node7_6 0 4.417545e-06
C6_8 node7_7 0 7.018853e-13
G6_8 node7_7 0 node7_7 0 4.410075e-06
C6_9 node7_8 0 6.973380e-13
G6_9 node7_8 0 node7_8 0 4.381504e-06
C6_10 node7_9 0 4.303249e-13
G6_10 node7_9 0 node7_9 0 2.703811e-06
CM6_1 node7_0 node7_1 -3.372270e-13
CM6_2 node7_0 node7_2 -4.333637e-14
CM6_3 node7_0 node7_3 -2.097687e-14
CM6_4 node7_0 node7_4 -1.177420e-14
CM6_5 node7_0 node7_5 -6.918544e-15
CM6_6 node7_0 node7_6 -4.146150e-15
CM6_7 node7_0 node7_7 -2.537949e-15
CM6_8 node7_0 node7_8 -1.643541e-15
CM6_9 node7_0 node7_9 -1.780983e-15
CM6_10 node7_1 node7_2 -3.044883e-13
CM6_11 node7_1 node7_3 -2.759806e-14
CM6_12 node7_1 node7_4 -1.220281e-14
CM6_13 node7_1 node7_5 -6.645893e-15
CM6_14 node7_1 node7_6 -3.879486e-15
CM6_15 node7_1 node7_7 -2.352696e-15
CM6_16 node7_1 node7_8 -1.518489e-15
CM6_17 node7_1 node7_9 -1.643380e-15
CM6_18 node7_2 node7_3 -3.019823e-13
CM6_19 node7_2 node7_4 -2.628447e-14
CM6_20 node7_2 node7_5 -1.143815e-14
CM6_21 node7_2 node7_6 -6.217217e-15
CM6_22 node7_2 node7_7 -3.678469e-15
CM6_23 node7_2 node7_8 -2.353400e-15
CM6_24 node7_2 node7_9 -2.538483e-15
CM6_25 node7_3 node7_4 -3.011554e-13
CM6_26 node7_3 node7_5 -2.592703e-14
CM6_27 node7_3 node7_6 -1.127554e-14
CM6_28 node7_3 node7_7 -6.213871e-15
CM6_29 node7_3 node7_8 -3.878491e-15
CM6_30 node7_3 node7_9 -4.144789e-15
CM6_31 node7_4 node7_5 -3.011387e-13
CM6_32 node7_4 node7_6 -2.590566e-14
CM6_33 node7_4 node7_7 -1.142857e-14
CM6_34 node7_4 node7_8 -6.642276e-15
CM6_35 node7_4 node7_9 -6.914501e-15
CM6_36 node7_5 node7_6 -3.012291e-13
CM6_37 node7_5 node7_7 -2.628136e-14
CM6_38 node7_5 node7_8 -1.220907e-14
CM6_39 node7_5 node7_9 -1.177964e-14
CM6_40 node7_6 node7_7 -3.018016e-13
CM6_41 node7_6 node7_8 -2.762580e-14
CM6_42 node7_6 node7_9 -2.099353e-14
CM6_43 node7_7 node7_8 -3.042640e-13
CM6_44 node7_7 node7_9 -4.332676e-14
CM6_45 node7_8 node7_9 -3.372029e-13
R7_1 node7_0 node7_0_mid 6.559697e-02
L7_1 node7_0_mid node8_0 1.324593e-01
R7_2 node7_1 node7_1_mid 6.559697e-02
L7_2 node7_1_mid node8_1 1.324593e-01
R7_3 node7_2 node7_2_mid 6.559697e-02
L7_3 node7_2_mid node8_2 1.324592e-01
R7_4 node7_3 node7_3_mid 6.559697e-02
L7_4 node7_3_mid node8_3 1.324592e-01
R7_5 node7_4 node7_4_mid 6.559697e-02
L7_5 node7_4_mid node8_4 1.324592e-01
R7_6 node7_5 node7_5_mid 6.559697e-02
L7_6 node7_5_mid node8_5 1.324591e-01
R7_7 node7_6 node7_6_mid 6.559697e-02
L7_7 node7_6_mid node8_6 1.324591e-01
R7_8 node7_7 node7_7_mid 6.559697e-02
L7_8 node7_7_mid node8_7 1.324591e-01
R7_9 node7_8 node7_8_mid 6.559697e-02
L7_9 node7_8_mid node8_8 1.324591e-01
R7_10 node7_9 node7_9_mid 6.559697e-02
L7_10 node7_9_mid node8_9 1.324591e-01
K7_1 L7_1 L7_2 1.000000e+00
K7_2 L7_1 L7_3 1.000000e+00
K7_3 L7_1 L7_4 1.000000e+00
K7_4 L7_1 L7_5 1.000000e+00
K7_5 L7_1 L7_6 9.999999e-01
K7_6 L7_1 L7_7 1.000000e+00
K7_7 L7_1 L7_8 9.999999e-01
K7_8 L7_1 L7_9 9.999999e-01
K7_9 L7_1 L7_10 9.999999e-01
K7_10 L7_2 L7_3 1.000000e+00
K7_11 L7_2 L7_4 1.000000e+00
K7_12 L7_2 L7_5 1.000000e+00
K7_13 L7_2 L7_6 9.999999e-01
K7_14 L7_2 L7_7 1.000000e+00
K7_15 L7_2 L7_8 9.999999e-01
K7_16 L7_2 L7_9 9.999999e-01
K7_17 L7_2 L7_10 9.999999e-01
K7_18 L7_3 L7_4 1.000000e+00
K7_19 L7_3 L7_5 1.000000e+00
K7_20 L7_3 L7_6 9.999999e-01
K7_21 L7_3 L7_7 9.999999e-01
K7_22 L7_3 L7_8 9.999999e-01
K7_23 L7_3 L7_9 9.999999e-01
K7_24 L7_3 L7_10 9.999998e-01
K7_25 L7_4 L7_5 1.000000e+00
K7_26 L7_4 L7_6 9.999999e-01
K7_27 L7_4 L7_7 1.000000e+00
K7_28 L7_4 L7_8 9.999999e-01
K7_29 L7_4 L7_9 9.999999e-01
K7_30 L7_4 L7_10 9.999999e-01
K7_31 L7_5 L7_6 9.999999e-01
K7_32 L7_5 L7_7 1.000000e+00
K7_33 L7_5 L7_8 9.999999e-01
K7_34 L7_5 L7_9 9.999999e-01
K7_35 L7_5 L7_10 9.999999e-01
K7_36 L7_6 L7_7 9.999999e-01
K7_37 L7_6 L7_8 1.000000e+00
K7_38 L7_6 L7_9 1.000000e+00
K7_39 L7_6 L7_10 9.999999e-01
K7_40 L7_7 L7_8 9.999999e-01
K7_41 L7_7 L7_9 9.999999e-01
K7_42 L7_7 L7_10 9.999999e-01
K7_43 L7_8 L7_9 1.000000e+00
K7_44 L7_8 L7_10 1.000000e+00
K7_45 L7_9 L7_10 1.000000e+00
C7_1 node8_0 0 4.303416e-13
G7_1 node8_0 0 node8_0 0 2.703916e-06
C7_2 node8_1 0 6.975560e-13
G7_2 node8_1 0 node8_1 0 4.382874e-06
C7_3 node8_2 0 7.023171e-13
G7_3 node8_2 0 node8_2 0 4.412789e-06
C7_4 node8_3 0 7.031524e-13
G7_4 node8_3 0 node8_3 0 4.418037e-06
C7_5 node8_4 0 7.034466e-13
G7_5 node8_4 0 node8_4 0 4.419885e-06
C7_6 node8_5 0 7.035676e-13
G7_6 node8_5 0 node8_5 0 4.420645e-06
C7_7 node8_6 0 7.030741e-13
G7_7 node8_6 0 node8_6 0 4.417545e-06
C7_8 node8_7 0 7.018853e-13
G7_8 node8_7 0 node8_7 0 4.410075e-06
C7_9 node8_8 0 6.973380e-13
G7_9 node8_8 0 node8_8 0 4.381504e-06
C7_10 node8_9 0 4.303249e-13
G7_10 node8_9 0 node8_9 0 2.703811e-06
CM7_1 node8_0 node8_1 -3.372270e-13
CM7_2 node8_0 node8_2 -4.333637e-14
CM7_3 node8_0 node8_3 -2.097687e-14
CM7_4 node8_0 node8_4 -1.177420e-14
CM7_5 node8_0 node8_5 -6.918544e-15
CM7_6 node8_0 node8_6 -4.146150e-15
CM7_7 node8_0 node8_7 -2.537949e-15
CM7_8 node8_0 node8_8 -1.643541e-15
CM7_9 node8_0 node8_9 -1.780983e-15
CM7_10 node8_1 node8_2 -3.044883e-13
CM7_11 node8_1 node8_3 -2.759806e-14
CM7_12 node8_1 node8_4 -1.220281e-14
CM7_13 node8_1 node8_5 -6.645893e-15
CM7_14 node8_1 node8_6 -3.879486e-15
CM7_15 node8_1 node8_7 -2.352696e-15
CM7_16 node8_1 node8_8 -1.518489e-15
CM7_17 node8_1 node8_9 -1.643380e-15
CM7_18 node8_2 node8_3 -3.019823e-13
CM7_19 node8_2 node8_4 -2.628447e-14
CM7_20 node8_2 node8_5 -1.143815e-14
CM7_21 node8_2 node8_6 -6.217217e-15
CM7_22 node8_2 node8_7 -3.678469e-15
CM7_23 node8_2 node8_8 -2.353400e-15
CM7_24 node8_2 node8_9 -2.538483e-15
CM7_25 node8_3 node8_4 -3.011554e-13
CM7_26 node8_3 node8_5 -2.592703e-14
CM7_27 node8_3 node8_6 -1.127554e-14
CM7_28 node8_3 node8_7 -6.213871e-15
CM7_29 node8_3 node8_8 -3.878491e-15
CM7_30 node8_3 node8_9 -4.144789e-15
CM7_31 node8_4 node8_5 -3.011387e-13
CM7_32 node8_4 node8_6 -2.590566e-14
CM7_33 node8_4 node8_7 -1.142857e-14
CM7_34 node8_4 node8_8 -6.642276e-15
CM7_35 node8_4 node8_9 -6.914501e-15
CM7_36 node8_5 node8_6 -3.012291e-13
CM7_37 node8_5 node8_7 -2.628136e-14
CM7_38 node8_5 node8_8 -1.220907e-14
CM7_39 node8_5 node8_9 -1.177964e-14
CM7_40 node8_6 node8_7 -3.018016e-13
CM7_41 node8_6 node8_8 -2.762580e-14
CM7_42 node8_6 node8_9 -2.099353e-14
CM7_43 node8_7 node8_8 -3.042640e-13
CM7_44 node8_7 node8_9 -4.332676e-14
CM7_45 node8_8 node8_9 -3.372029e-13
R8_1 node8_0 node8_0_mid 6.559697e-02
L8_1 node8_0_mid node9_0 1.324593e-01
R8_2 node8_1 node8_1_mid 6.559697e-02
L8_2 node8_1_mid node9_1 1.324593e-01
R8_3 node8_2 node8_2_mid 6.559697e-02
L8_3 node8_2_mid node9_2 1.324592e-01
R8_4 node8_3 node8_3_mid 6.559697e-02
L8_4 node8_3_mid node9_3 1.324592e-01
R8_5 node8_4 node8_4_mid 6.559697e-02
L8_5 node8_4_mid node9_4 1.324592e-01
R8_6 node8_5 node8_5_mid 6.559697e-02
L8_6 node8_5_mid node9_5 1.324591e-01
R8_7 node8_6 node8_6_mid 6.559697e-02
L8_7 node8_6_mid node9_6 1.324591e-01
R8_8 node8_7 node8_7_mid 6.559697e-02
L8_8 node8_7_mid node9_7 1.324591e-01
R8_9 node8_8 node8_8_mid 6.559697e-02
L8_9 node8_8_mid node9_8 1.324591e-01
R8_10 node8_9 node8_9_mid 6.559697e-02
L8_10 node8_9_mid node9_9 1.324591e-01
K8_1 L8_1 L8_2 1.000000e+00
K8_2 L8_1 L8_3 1.000000e+00
K8_3 L8_1 L8_4 1.000000e+00
K8_4 L8_1 L8_5 1.000000e+00
K8_5 L8_1 L8_6 9.999999e-01
K8_6 L8_1 L8_7 1.000000e+00
K8_7 L8_1 L8_8 9.999999e-01
K8_8 L8_1 L8_9 9.999999e-01
K8_9 L8_1 L8_10 9.999999e-01
K8_10 L8_2 L8_3 1.000000e+00
K8_11 L8_2 L8_4 1.000000e+00
K8_12 L8_2 L8_5 1.000000e+00
K8_13 L8_2 L8_6 9.999999e-01
K8_14 L8_2 L8_7 1.000000e+00
K8_15 L8_2 L8_8 9.999999e-01
K8_16 L8_2 L8_9 9.999999e-01
K8_17 L8_2 L8_10 9.999999e-01
K8_18 L8_3 L8_4 1.000000e+00
K8_19 L8_3 L8_5 1.000000e+00
K8_20 L8_3 L8_6 9.999999e-01
K8_21 L8_3 L8_7 9.999999e-01
K8_22 L8_3 L8_8 9.999999e-01
K8_23 L8_3 L8_9 9.999999e-01
K8_24 L8_3 L8_10 9.999998e-01
K8_25 L8_4 L8_5 1.000000e+00
K8_26 L8_4 L8_6 9.999999e-01
K8_27 L8_4 L8_7 1.000000e+00
K8_28 L8_4 L8_8 9.999999e-01
K8_29 L8_4 L8_9 9.999999e-01
K8_30 L8_4 L8_10 9.999999e-01
K8_31 L8_5 L8_6 9.999999e-01
K8_32 L8_5 L8_7 1.000000e+00
K8_33 L8_5 L8_8 9.999999e-01
K8_34 L8_5 L8_9 9.999999e-01
K8_35 L8_5 L8_10 9.999999e-01
K8_36 L8_6 L8_7 9.999999e-01
K8_37 L8_6 L8_8 1.000000e+00
K8_38 L8_6 L8_9 1.000000e+00
K8_39 L8_6 L8_10 9.999999e-01
K8_40 L8_7 L8_8 9.999999e-01
K8_41 L8_7 L8_9 9.999999e-01
K8_42 L8_7 L8_10 9.999999e-01
K8_43 L8_8 L8_9 1.000000e+00
K8_44 L8_8 L8_10 1.000000e+00
K8_45 L8_9 L8_10 1.000000e+00
C8_1 node9_0 0 4.303416e-13
G8_1 node9_0 0 node9_0 0 2.703916e-06
C8_2 node9_1 0 6.975560e-13
G8_2 node9_1 0 node9_1 0 4.382874e-06
C8_3 node9_2 0 7.023171e-13
G8_3 node9_2 0 node9_2 0 4.412789e-06
C8_4 node9_3 0 7.031524e-13
G8_4 node9_3 0 node9_3 0 4.418037e-06
C8_5 node9_4 0 7.034466e-13
G8_5 node9_4 0 node9_4 0 4.419885e-06
C8_6 node9_5 0 7.035676e-13
G8_6 node9_5 0 node9_5 0 4.420645e-06
C8_7 node9_6 0 7.030741e-13
G8_7 node9_6 0 node9_6 0 4.417545e-06
C8_8 node9_7 0 7.018853e-13
G8_8 node9_7 0 node9_7 0 4.410075e-06
C8_9 node9_8 0 6.973380e-13
G8_9 node9_8 0 node9_8 0 4.381504e-06
C8_10 node9_9 0 4.303249e-13
G8_10 node9_9 0 node9_9 0 2.703811e-06
CM8_1 node9_0 node9_1 -3.372270e-13
CM8_2 node9_0 node9_2 -4.333637e-14
CM8_3 node9_0 node9_3 -2.097687e-14
CM8_4 node9_0 node9_4 -1.177420e-14
CM8_5 node9_0 node9_5 -6.918544e-15
CM8_6 node9_0 node9_6 -4.146150e-15
CM8_7 node9_0 node9_7 -2.537949e-15
CM8_8 node9_0 node9_8 -1.643541e-15
CM8_9 node9_0 node9_9 -1.780983e-15
CM8_10 node9_1 node9_2 -3.044883e-13
CM8_11 node9_1 node9_3 -2.759806e-14
CM8_12 node9_1 node9_4 -1.220281e-14
CM8_13 node9_1 node9_5 -6.645893e-15
CM8_14 node9_1 node9_6 -3.879486e-15
CM8_15 node9_1 node9_7 -2.352696e-15
CM8_16 node9_1 node9_8 -1.518489e-15
CM8_17 node9_1 node9_9 -1.643380e-15
CM8_18 node9_2 node9_3 -3.019823e-13
CM8_19 node9_2 node9_4 -2.628447e-14
CM8_20 node9_2 node9_5 -1.143815e-14
CM8_21 node9_2 node9_6 -6.217217e-15
CM8_22 node9_2 node9_7 -3.678469e-15
CM8_23 node9_2 node9_8 -2.353400e-15
CM8_24 node9_2 node9_9 -2.538483e-15
CM8_25 node9_3 node9_4 -3.011554e-13
CM8_26 node9_3 node9_5 -2.592703e-14
CM8_27 node9_3 node9_6 -1.127554e-14
CM8_28 node9_3 node9_7 -6.213871e-15
CM8_29 node9_3 node9_8 -3.878491e-15
CM8_30 node9_3 node9_9 -4.144789e-15
CM8_31 node9_4 node9_5 -3.011387e-13
CM8_32 node9_4 node9_6 -2.590566e-14
CM8_33 node9_4 node9_7 -1.142857e-14
CM8_34 node9_4 node9_8 -6.642276e-15
CM8_35 node9_4 node9_9 -6.914501e-15
CM8_36 node9_5 node9_6 -3.012291e-13
CM8_37 node9_5 node9_7 -2.628136e-14
CM8_38 node9_5 node9_8 -1.220907e-14
CM8_39 node9_5 node9_9 -1.177964e-14
CM8_40 node9_6 node9_7 -3.018016e-13
CM8_41 node9_6 node9_8 -2.762580e-14
CM8_42 node9_6 node9_9 -2.099353e-14
CM8_43 node9_7 node9_8 -3.042640e-13
CM8_44 node9_7 node9_9 -4.332676e-14
CM8_45 node9_8 node9_9 -3.372029e-13
R9_1 node9_0 node9_0_mid 6.559697e-02
L9_1 node9_0_mid node10_0 1.324593e-01
R9_2 node9_1 node9_1_mid 6.559697e-02
L9_2 node9_1_mid node10_1 1.324593e-01
R9_3 node9_2 node9_2_mid 6.559697e-02
L9_3 node9_2_mid node10_2 1.324592e-01
R9_4 node9_3 node9_3_mid 6.559697e-02
L9_4 node9_3_mid node10_3 1.324592e-01
R9_5 node9_4 node9_4_mid 6.559697e-02
L9_5 node9_4_mid node10_4 1.324592e-01
R9_6 node9_5 node9_5_mid 6.559697e-02
L9_6 node9_5_mid node10_5 1.324591e-01
R9_7 node9_6 node9_6_mid 6.559697e-02
L9_7 node9_6_mid node10_6 1.324591e-01
R9_8 node9_7 node9_7_mid 6.559697e-02
L9_8 node9_7_mid node10_7 1.324591e-01
R9_9 node9_8 node9_8_mid 6.559697e-02
L9_9 node9_8_mid node10_8 1.324591e-01
R9_10 node9_9 node9_9_mid 6.559697e-02
L9_10 node9_9_mid node10_9 1.324591e-01
K9_1 L9_1 L9_2 1.000000e+00
K9_2 L9_1 L9_3 1.000000e+00
K9_3 L9_1 L9_4 1.000000e+00
K9_4 L9_1 L9_5 1.000000e+00
K9_5 L9_1 L9_6 9.999999e-01
K9_6 L9_1 L9_7 1.000000e+00
K9_7 L9_1 L9_8 9.999999e-01
K9_8 L9_1 L9_9 9.999999e-01
K9_9 L9_1 L9_10 9.999999e-01
K9_10 L9_2 L9_3 1.000000e+00
K9_11 L9_2 L9_4 1.000000e+00
K9_12 L9_2 L9_5 1.000000e+00
K9_13 L9_2 L9_6 9.999999e-01
K9_14 L9_2 L9_7 1.000000e+00
K9_15 L9_2 L9_8 9.999999e-01
K9_16 L9_2 L9_9 9.999999e-01
K9_17 L9_2 L9_10 9.999999e-01
K9_18 L9_3 L9_4 1.000000e+00
K9_19 L9_3 L9_5 1.000000e+00
K9_20 L9_3 L9_6 9.999999e-01
K9_21 L9_3 L9_7 9.999999e-01
K9_22 L9_3 L9_8 9.999999e-01
K9_23 L9_3 L9_9 9.999999e-01
K9_24 L9_3 L9_10 9.999998e-01
K9_25 L9_4 L9_5 1.000000e+00
K9_26 L9_4 L9_6 9.999999e-01
K9_27 L9_4 L9_7 1.000000e+00
K9_28 L9_4 L9_8 9.999999e-01
K9_29 L9_4 L9_9 9.999999e-01
K9_30 L9_4 L9_10 9.999999e-01
K9_31 L9_5 L9_6 9.999999e-01
K9_32 L9_5 L9_7 1.000000e+00
K9_33 L9_5 L9_8 9.999999e-01
K9_34 L9_5 L9_9 9.999999e-01
K9_35 L9_5 L9_10 9.999999e-01
K9_36 L9_6 L9_7 9.999999e-01
K9_37 L9_6 L9_8 1.000000e+00
K9_38 L9_6 L9_9 1.000000e+00
K9_39 L9_6 L9_10 9.999999e-01
K9_40 L9_7 L9_8 9.999999e-01
K9_41 L9_7 L9_9 9.999999e-01
K9_42 L9_7 L9_10 9.999999e-01
K9_43 L9_8 L9_9 1.000000e+00
K9_44 L9_8 L9_10 1.000000e+00
K9_45 L9_9 L9_10 1.000000e+00
C9_1 node10_0 0 4.303416e-13
G9_1 node10_0 0 node10_0 0 2.703916e-06
C9_2 node10_1 0 6.975560e-13
G9_2 node10_1 0 node10_1 0 4.382874e-06
C9_3 node10_2 0 7.023171e-13
G9_3 node10_2 0 node10_2 0 4.412789e-06
C9_4 node10_3 0 7.031524e-13
G9_4 node10_3 0 node10_3 0 4.418037e-06
C9_5 node10_4 0 7.034466e-13
G9_5 node10_4 0 node10_4 0 4.419885e-06
C9_6 node10_5 0 7.035676e-13
G9_6 node10_5 0 node10_5 0 4.420645e-06
C9_7 node10_6 0 7.030741e-13
G9_7 node10_6 0 node10_6 0 4.417545e-06
C9_8 node10_7 0 7.018853e-13
G9_8 node10_7 0 node10_7 0 4.410075e-06
C9_9 node10_8 0 6.973380e-13
G9_9 node10_8 0 node10_8 0 4.381504e-06
C9_10 node10_9 0 4.303249e-13
G9_10 node10_9 0 node10_9 0 2.703811e-06
CM9_1 node10_0 node10_1 -3.372270e-13
CM9_2 node10_0 node10_2 -4.333637e-14
CM9_3 node10_0 node10_3 -2.097687e-14
CM9_4 node10_0 node10_4 -1.177420e-14
CM9_5 node10_0 node10_5 -6.918544e-15
CM9_6 node10_0 node10_6 -4.146150e-15
CM9_7 node10_0 node10_7 -2.537949e-15
CM9_8 node10_0 node10_8 -1.643541e-15
CM9_9 node10_0 node10_9 -1.780983e-15
CM9_10 node10_1 node10_2 -3.044883e-13
CM9_11 node10_1 node10_3 -2.759806e-14
CM9_12 node10_1 node10_4 -1.220281e-14
CM9_13 node10_1 node10_5 -6.645893e-15
CM9_14 node10_1 node10_6 -3.879486e-15
CM9_15 node10_1 node10_7 -2.352696e-15
CM9_16 node10_1 node10_8 -1.518489e-15
CM9_17 node10_1 node10_9 -1.643380e-15
CM9_18 node10_2 node10_3 -3.019823e-13
CM9_19 node10_2 node10_4 -2.628447e-14
CM9_20 node10_2 node10_5 -1.143815e-14
CM9_21 node10_2 node10_6 -6.217217e-15
CM9_22 node10_2 node10_7 -3.678469e-15
CM9_23 node10_2 node10_8 -2.353400e-15
CM9_24 node10_2 node10_9 -2.538483e-15
CM9_25 node10_3 node10_4 -3.011554e-13
CM9_26 node10_3 node10_5 -2.592703e-14
CM9_27 node10_3 node10_6 -1.127554e-14
CM9_28 node10_3 node10_7 -6.213871e-15
CM9_29 node10_3 node10_8 -3.878491e-15
CM9_30 node10_3 node10_9 -4.144789e-15
CM9_31 node10_4 node10_5 -3.011387e-13
CM9_32 node10_4 node10_6 -2.590566e-14
CM9_33 node10_4 node10_7 -1.142857e-14
CM9_34 node10_4 node10_8 -6.642276e-15
CM9_35 node10_4 node10_9 -6.914501e-15
CM9_36 node10_5 node10_6 -3.012291e-13
CM9_37 node10_5 node10_7 -2.628136e-14
CM9_38 node10_5 node10_8 -1.220907e-14
CM9_39 node10_5 node10_9 -1.177964e-14
CM9_40 node10_6 node10_7 -3.018016e-13
CM9_41 node10_6 node10_8 -2.762580e-14
CM9_42 node10_6 node10_9 -2.099353e-14
CM9_43 node10_7 node10_8 -3.042640e-13
CM9_44 node10_7 node10_9 -4.332676e-14
CM9_45 node10_8 node10_9 -3.372029e-13
R10_1 node10_0 node10_0_mid 6.559697e-02
L10_1 node10_0_mid node11_0 1.324593e-01
R10_2 node10_1 node10_1_mid 6.559697e-02
L10_2 node10_1_mid node11_1 1.324593e-01
R10_3 node10_2 node10_2_mid 6.559697e-02
L10_3 node10_2_mid node11_2 1.324592e-01
R10_4 node10_3 node10_3_mid 6.559697e-02
L10_4 node10_3_mid node11_3 1.324592e-01
R10_5 node10_4 node10_4_mid 6.559697e-02
L10_5 node10_4_mid node11_4 1.324592e-01
R10_6 node10_5 node10_5_mid 6.559697e-02
L10_6 node10_5_mid node11_5 1.324591e-01
R10_7 node10_6 node10_6_mid 6.559697e-02
L10_7 node10_6_mid node11_6 1.324591e-01
R10_8 node10_7 node10_7_mid 6.559697e-02
L10_8 node10_7_mid node11_7 1.324591e-01
R10_9 node10_8 node10_8_mid 6.559697e-02
L10_9 node10_8_mid node11_8 1.324591e-01
R10_10 node10_9 node10_9_mid 6.559697e-02
L10_10 node10_9_mid node11_9 1.324591e-01
K10_1 L10_1 L10_2 1.000000e+00
K10_2 L10_1 L10_3 1.000000e+00
K10_3 L10_1 L10_4 1.000000e+00
K10_4 L10_1 L10_5 1.000000e+00
K10_5 L10_1 L10_6 9.999999e-01
K10_6 L10_1 L10_7 1.000000e+00
K10_7 L10_1 L10_8 9.999999e-01
K10_8 L10_1 L10_9 9.999999e-01
K10_9 L10_1 L10_10 9.999999e-01
K10_10 L10_2 L10_3 1.000000e+00
K10_11 L10_2 L10_4 1.000000e+00
K10_12 L10_2 L10_5 1.000000e+00
K10_13 L10_2 L10_6 9.999999e-01
K10_14 L10_2 L10_7 1.000000e+00
K10_15 L10_2 L10_8 9.999999e-01
K10_16 L10_2 L10_9 9.999999e-01
K10_17 L10_2 L10_10 9.999999e-01
K10_18 L10_3 L10_4 1.000000e+00
K10_19 L10_3 L10_5 1.000000e+00
K10_20 L10_3 L10_6 9.999999e-01
K10_21 L10_3 L10_7 9.999999e-01
K10_22 L10_3 L10_8 9.999999e-01
K10_23 L10_3 L10_9 9.999999e-01
K10_24 L10_3 L10_10 9.999998e-01
K10_25 L10_4 L10_5 1.000000e+00
K10_26 L10_4 L10_6 9.999999e-01
K10_27 L10_4 L10_7 1.000000e+00
K10_28 L10_4 L10_8 9.999999e-01
K10_29 L10_4 L10_9 9.999999e-01
K10_30 L10_4 L10_10 9.999999e-01
K10_31 L10_5 L10_6 9.999999e-01
K10_32 L10_5 L10_7 1.000000e+00
K10_33 L10_5 L10_8 9.999999e-01
K10_34 L10_5 L10_9 9.999999e-01
K10_35 L10_5 L10_10 9.999999e-01
K10_36 L10_6 L10_7 9.999999e-01
K10_37 L10_6 L10_8 1.000000e+00
K10_38 L10_6 L10_9 1.000000e+00
K10_39 L10_6 L10_10 9.999999e-01
K10_40 L10_7 L10_8 9.999999e-01
K10_41 L10_7 L10_9 9.999999e-01
K10_42 L10_7 L10_10 9.999999e-01
K10_43 L10_8 L10_9 1.000000e+00
K10_44 L10_8 L10_10 1.000000e+00
K10_45 L10_9 L10_10 1.000000e+00
C10_1 node11_0 0 4.303416e-13
G10_1 node11_0 0 node11_0 0 2.703916e-06
C10_2 node11_1 0 6.975560e-13
G10_2 node11_1 0 node11_1 0 4.382874e-06
C10_3 node11_2 0 7.023171e-13
G10_3 node11_2 0 node11_2 0 4.412789e-06
C10_4 node11_3 0 7.031524e-13
G10_4 node11_3 0 node11_3 0 4.418037e-06
C10_5 node11_4 0 7.034466e-13
G10_5 node11_4 0 node11_4 0 4.419885e-06
C10_6 node11_5 0 7.035676e-13
G10_6 node11_5 0 node11_5 0 4.420645e-06
C10_7 node11_6 0 7.030741e-13
G10_7 node11_6 0 node11_6 0 4.417545e-06
C10_8 node11_7 0 7.018853e-13
G10_8 node11_7 0 node11_7 0 4.410075e-06
C10_9 node11_8 0 6.973380e-13
G10_9 node11_8 0 node11_8 0 4.381504e-06
C10_10 node11_9 0 4.303249e-13
G10_10 node11_9 0 node11_9 0 2.703811e-06
CM10_1 node11_0 node11_1 -3.372270e-13
CM10_2 node11_0 node11_2 -4.333637e-14
CM10_3 node11_0 node11_3 -2.097687e-14
CM10_4 node11_0 node11_4 -1.177420e-14
CM10_5 node11_0 node11_5 -6.918544e-15
CM10_6 node11_0 node11_6 -4.146150e-15
CM10_7 node11_0 node11_7 -2.537949e-15
CM10_8 node11_0 node11_8 -1.643541e-15
CM10_9 node11_0 node11_9 -1.780983e-15
CM10_10 node11_1 node11_2 -3.044883e-13
CM10_11 node11_1 node11_3 -2.759806e-14
CM10_12 node11_1 node11_4 -1.220281e-14
CM10_13 node11_1 node11_5 -6.645893e-15
CM10_14 node11_1 node11_6 -3.879486e-15
CM10_15 node11_1 node11_7 -2.352696e-15
CM10_16 node11_1 node11_8 -1.518489e-15
CM10_17 node11_1 node11_9 -1.643380e-15
CM10_18 node11_2 node11_3 -3.019823e-13
CM10_19 node11_2 node11_4 -2.628447e-14
CM10_20 node11_2 node11_5 -1.143815e-14
CM10_21 node11_2 node11_6 -6.217217e-15
CM10_22 node11_2 node11_7 -3.678469e-15
CM10_23 node11_2 node11_8 -2.353400e-15
CM10_24 node11_2 node11_9 -2.538483e-15
CM10_25 node11_3 node11_4 -3.011554e-13
CM10_26 node11_3 node11_5 -2.592703e-14
CM10_27 node11_3 node11_6 -1.127554e-14
CM10_28 node11_3 node11_7 -6.213871e-15
CM10_29 node11_3 node11_8 -3.878491e-15
CM10_30 node11_3 node11_9 -4.144789e-15
CM10_31 node11_4 node11_5 -3.011387e-13
CM10_32 node11_4 node11_6 -2.590566e-14
CM10_33 node11_4 node11_7 -1.142857e-14
CM10_34 node11_4 node11_8 -6.642276e-15
CM10_35 node11_4 node11_9 -6.914501e-15
CM10_36 node11_5 node11_6 -3.012291e-13
CM10_37 node11_5 node11_7 -2.628136e-14
CM10_38 node11_5 node11_8 -1.220907e-14
CM10_39 node11_5 node11_9 -1.177964e-14
CM10_40 node11_6 node11_7 -3.018016e-13
CM10_41 node11_6 node11_8 -2.762580e-14
CM10_42 node11_6 node11_9 -2.099353e-14
CM10_43 node11_7 node11_8 -3.042640e-13
CM10_44 node11_7 node11_9 -4.332676e-14
CM10_45 node11_8 node11_9 -3.372029e-13
R11_1 node11_0 node11_0_mid 6.559697e-02
L11_1 node11_0_mid node12_0 1.324593e-01
R11_2 node11_1 node11_1_mid 6.559697e-02
L11_2 node11_1_mid node12_1 1.324593e-01
R11_3 node11_2 node11_2_mid 6.559697e-02
L11_3 node11_2_mid node12_2 1.324592e-01
R11_4 node11_3 node11_3_mid 6.559697e-02
L11_4 node11_3_mid node12_3 1.324592e-01
R11_5 node11_4 node11_4_mid 6.559697e-02
L11_5 node11_4_mid node12_4 1.324592e-01
R11_6 node11_5 node11_5_mid 6.559697e-02
L11_6 node11_5_mid node12_5 1.324591e-01
R11_7 node11_6 node11_6_mid 6.559697e-02
L11_7 node11_6_mid node12_6 1.324591e-01
R11_8 node11_7 node11_7_mid 6.559697e-02
L11_8 node11_7_mid node12_7 1.324591e-01
R11_9 node11_8 node11_8_mid 6.559697e-02
L11_9 node11_8_mid node12_8 1.324591e-01
R11_10 node11_9 node11_9_mid 6.559697e-02
L11_10 node11_9_mid node12_9 1.324591e-01
K11_1 L11_1 L11_2 1.000000e+00
K11_2 L11_1 L11_3 1.000000e+00
K11_3 L11_1 L11_4 1.000000e+00
K11_4 L11_1 L11_5 1.000000e+00
K11_5 L11_1 L11_6 9.999999e-01
K11_6 L11_1 L11_7 1.000000e+00
K11_7 L11_1 L11_8 9.999999e-01
K11_8 L11_1 L11_9 9.999999e-01
K11_9 L11_1 L11_10 9.999999e-01
K11_10 L11_2 L11_3 1.000000e+00
K11_11 L11_2 L11_4 1.000000e+00
K11_12 L11_2 L11_5 1.000000e+00
K11_13 L11_2 L11_6 9.999999e-01
K11_14 L11_2 L11_7 1.000000e+00
K11_15 L11_2 L11_8 9.999999e-01
K11_16 L11_2 L11_9 9.999999e-01
K11_17 L11_2 L11_10 9.999999e-01
K11_18 L11_3 L11_4 1.000000e+00
K11_19 L11_3 L11_5 1.000000e+00
K11_20 L11_3 L11_6 9.999999e-01
K11_21 L11_3 L11_7 9.999999e-01
K11_22 L11_3 L11_8 9.999999e-01
K11_23 L11_3 L11_9 9.999999e-01
K11_24 L11_3 L11_10 9.999998e-01
K11_25 L11_4 L11_5 1.000000e+00
K11_26 L11_4 L11_6 9.999999e-01
K11_27 L11_4 L11_7 1.000000e+00
K11_28 L11_4 L11_8 9.999999e-01
K11_29 L11_4 L11_9 9.999999e-01
K11_30 L11_4 L11_10 9.999999e-01
K11_31 L11_5 L11_6 9.999999e-01
K11_32 L11_5 L11_7 1.000000e+00
K11_33 L11_5 L11_8 9.999999e-01
K11_34 L11_5 L11_9 9.999999e-01
K11_35 L11_5 L11_10 9.999999e-01
K11_36 L11_6 L11_7 9.999999e-01
K11_37 L11_6 L11_8 1.000000e+00
K11_38 L11_6 L11_9 1.000000e+00
K11_39 L11_6 L11_10 9.999999e-01
K11_40 L11_7 L11_8 9.999999e-01
K11_41 L11_7 L11_9 9.999999e-01
K11_42 L11_7 L11_10 9.999999e-01
K11_43 L11_8 L11_9 1.000000e+00
K11_44 L11_8 L11_10 1.000000e+00
K11_45 L11_9 L11_10 1.000000e+00
C11_1 node12_0 0 4.303416e-13
G11_1 node12_0 0 node12_0 0 2.703916e-06
C11_2 node12_1 0 6.975560e-13
G11_2 node12_1 0 node12_1 0 4.382874e-06
C11_3 node12_2 0 7.023171e-13
G11_3 node12_2 0 node12_2 0 4.412789e-06
C11_4 node12_3 0 7.031524e-13
G11_4 node12_3 0 node12_3 0 4.418037e-06
C11_5 node12_4 0 7.034466e-13
G11_5 node12_4 0 node12_4 0 4.419885e-06
C11_6 node12_5 0 7.035676e-13
G11_6 node12_5 0 node12_5 0 4.420645e-06
C11_7 node12_6 0 7.030741e-13
G11_7 node12_6 0 node12_6 0 4.417545e-06
C11_8 node12_7 0 7.018853e-13
G11_8 node12_7 0 node12_7 0 4.410075e-06
C11_9 node12_8 0 6.973380e-13
G11_9 node12_8 0 node12_8 0 4.381504e-06
C11_10 node12_9 0 4.303249e-13
G11_10 node12_9 0 node12_9 0 2.703811e-06
CM11_1 node12_0 node12_1 -3.372270e-13
CM11_2 node12_0 node12_2 -4.333637e-14
CM11_3 node12_0 node12_3 -2.097687e-14
CM11_4 node12_0 node12_4 -1.177420e-14
CM11_5 node12_0 node12_5 -6.918544e-15
CM11_6 node12_0 node12_6 -4.146150e-15
CM11_7 node12_0 node12_7 -2.537949e-15
CM11_8 node12_0 node12_8 -1.643541e-15
CM11_9 node12_0 node12_9 -1.780983e-15
CM11_10 node12_1 node12_2 -3.044883e-13
CM11_11 node12_1 node12_3 -2.759806e-14
CM11_12 node12_1 node12_4 -1.220281e-14
CM11_13 node12_1 node12_5 -6.645893e-15
CM11_14 node12_1 node12_6 -3.879486e-15
CM11_15 node12_1 node12_7 -2.352696e-15
CM11_16 node12_1 node12_8 -1.518489e-15
CM11_17 node12_1 node12_9 -1.643380e-15
CM11_18 node12_2 node12_3 -3.019823e-13
CM11_19 node12_2 node12_4 -2.628447e-14
CM11_20 node12_2 node12_5 -1.143815e-14
CM11_21 node12_2 node12_6 -6.217217e-15
CM11_22 node12_2 node12_7 -3.678469e-15
CM11_23 node12_2 node12_8 -2.353400e-15
CM11_24 node12_2 node12_9 -2.538483e-15
CM11_25 node12_3 node12_4 -3.011554e-13
CM11_26 node12_3 node12_5 -2.592703e-14
CM11_27 node12_3 node12_6 -1.127554e-14
CM11_28 node12_3 node12_7 -6.213871e-15
CM11_29 node12_3 node12_8 -3.878491e-15
CM11_30 node12_3 node12_9 -4.144789e-15
CM11_31 node12_4 node12_5 -3.011387e-13
CM11_32 node12_4 node12_6 -2.590566e-14
CM11_33 node12_4 node12_7 -1.142857e-14
CM11_34 node12_4 node12_8 -6.642276e-15
CM11_35 node12_4 node12_9 -6.914501e-15
CM11_36 node12_5 node12_6 -3.012291e-13
CM11_37 node12_5 node12_7 -2.628136e-14
CM11_38 node12_5 node12_8 -1.220907e-14
CM11_39 node12_5 node12_9 -1.177964e-14
CM11_40 node12_6 node12_7 -3.018016e-13
CM11_41 node12_6 node12_8 -2.762580e-14
CM11_42 node12_6 node12_9 -2.099353e-14
CM11_43 node12_7 node12_8 -3.042640e-13
CM11_44 node12_7 node12_9 -4.332676e-14
CM11_45 node12_8 node12_9 -3.372029e-13
R12_1 node12_0 node12_0_mid 6.559697e-02
L12_1 node12_0_mid node13_0 1.324593e-01
R12_2 node12_1 node12_1_mid 6.559697e-02
L12_2 node12_1_mid node13_1 1.324593e-01
R12_3 node12_2 node12_2_mid 6.559697e-02
L12_3 node12_2_mid node13_2 1.324592e-01
R12_4 node12_3 node12_3_mid 6.559697e-02
L12_4 node12_3_mid node13_3 1.324592e-01
R12_5 node12_4 node12_4_mid 6.559697e-02
L12_5 node12_4_mid node13_4 1.324592e-01
R12_6 node12_5 node12_5_mid 6.559697e-02
L12_6 node12_5_mid node13_5 1.324591e-01
R12_7 node12_6 node12_6_mid 6.559697e-02
L12_7 node12_6_mid node13_6 1.324591e-01
R12_8 node12_7 node12_7_mid 6.559697e-02
L12_8 node12_7_mid node13_7 1.324591e-01
R12_9 node12_8 node12_8_mid 6.559697e-02
L12_9 node12_8_mid node13_8 1.324591e-01
R12_10 node12_9 node12_9_mid 6.559697e-02
L12_10 node12_9_mid node13_9 1.324591e-01
K12_1 L12_1 L12_2 1.000000e+00
K12_2 L12_1 L12_3 1.000000e+00
K12_3 L12_1 L12_4 1.000000e+00
K12_4 L12_1 L12_5 1.000000e+00
K12_5 L12_1 L12_6 9.999999e-01
K12_6 L12_1 L12_7 1.000000e+00
K12_7 L12_1 L12_8 9.999999e-01
K12_8 L12_1 L12_9 9.999999e-01
K12_9 L12_1 L12_10 9.999999e-01
K12_10 L12_2 L12_3 1.000000e+00
K12_11 L12_2 L12_4 1.000000e+00
K12_12 L12_2 L12_5 1.000000e+00
K12_13 L12_2 L12_6 9.999999e-01
K12_14 L12_2 L12_7 1.000000e+00
K12_15 L12_2 L12_8 9.999999e-01
K12_16 L12_2 L12_9 9.999999e-01
K12_17 L12_2 L12_10 9.999999e-01
K12_18 L12_3 L12_4 1.000000e+00
K12_19 L12_3 L12_5 1.000000e+00
K12_20 L12_3 L12_6 9.999999e-01
K12_21 L12_3 L12_7 9.999999e-01
K12_22 L12_3 L12_8 9.999999e-01
K12_23 L12_3 L12_9 9.999999e-01
K12_24 L12_3 L12_10 9.999998e-01
K12_25 L12_4 L12_5 1.000000e+00
K12_26 L12_4 L12_6 9.999999e-01
K12_27 L12_4 L12_7 1.000000e+00
K12_28 L12_4 L12_8 9.999999e-01
K12_29 L12_4 L12_9 9.999999e-01
K12_30 L12_4 L12_10 9.999999e-01
K12_31 L12_5 L12_6 9.999999e-01
K12_32 L12_5 L12_7 1.000000e+00
K12_33 L12_5 L12_8 9.999999e-01
K12_34 L12_5 L12_9 9.999999e-01
K12_35 L12_5 L12_10 9.999999e-01
K12_36 L12_6 L12_7 9.999999e-01
K12_37 L12_6 L12_8 1.000000e+00
K12_38 L12_6 L12_9 1.000000e+00
K12_39 L12_6 L12_10 9.999999e-01
K12_40 L12_7 L12_8 9.999999e-01
K12_41 L12_7 L12_9 9.999999e-01
K12_42 L12_7 L12_10 9.999999e-01
K12_43 L12_8 L12_9 1.000000e+00
K12_44 L12_8 L12_10 1.000000e+00
K12_45 L12_9 L12_10 1.000000e+00
C12_1 node13_0 0 4.303416e-13
G12_1 node13_0 0 node13_0 0 2.703916e-06
C12_2 node13_1 0 6.975560e-13
G12_2 node13_1 0 node13_1 0 4.382874e-06
C12_3 node13_2 0 7.023171e-13
G12_3 node13_2 0 node13_2 0 4.412789e-06
C12_4 node13_3 0 7.031524e-13
G12_4 node13_3 0 node13_3 0 4.418037e-06
C12_5 node13_4 0 7.034466e-13
G12_5 node13_4 0 node13_4 0 4.419885e-06
C12_6 node13_5 0 7.035676e-13
G12_6 node13_5 0 node13_5 0 4.420645e-06
C12_7 node13_6 0 7.030741e-13
G12_7 node13_6 0 node13_6 0 4.417545e-06
C12_8 node13_7 0 7.018853e-13
G12_8 node13_7 0 node13_7 0 4.410075e-06
C12_9 node13_8 0 6.973380e-13
G12_9 node13_8 0 node13_8 0 4.381504e-06
C12_10 node13_9 0 4.303249e-13
G12_10 node13_9 0 node13_9 0 2.703811e-06
CM12_1 node13_0 node13_1 -3.372270e-13
CM12_2 node13_0 node13_2 -4.333637e-14
CM12_3 node13_0 node13_3 -2.097687e-14
CM12_4 node13_0 node13_4 -1.177420e-14
CM12_5 node13_0 node13_5 -6.918544e-15
CM12_6 node13_0 node13_6 -4.146150e-15
CM12_7 node13_0 node13_7 -2.537949e-15
CM12_8 node13_0 node13_8 -1.643541e-15
CM12_9 node13_0 node13_9 -1.780983e-15
CM12_10 node13_1 node13_2 -3.044883e-13
CM12_11 node13_1 node13_3 -2.759806e-14
CM12_12 node13_1 node13_4 -1.220281e-14
CM12_13 node13_1 node13_5 -6.645893e-15
CM12_14 node13_1 node13_6 -3.879486e-15
CM12_15 node13_1 node13_7 -2.352696e-15
CM12_16 node13_1 node13_8 -1.518489e-15
CM12_17 node13_1 node13_9 -1.643380e-15
CM12_18 node13_2 node13_3 -3.019823e-13
CM12_19 node13_2 node13_4 -2.628447e-14
CM12_20 node13_2 node13_5 -1.143815e-14
CM12_21 node13_2 node13_6 -6.217217e-15
CM12_22 node13_2 node13_7 -3.678469e-15
CM12_23 node13_2 node13_8 -2.353400e-15
CM12_24 node13_2 node13_9 -2.538483e-15
CM12_25 node13_3 node13_4 -3.011554e-13
CM12_26 node13_3 node13_5 -2.592703e-14
CM12_27 node13_3 node13_6 -1.127554e-14
CM12_28 node13_3 node13_7 -6.213871e-15
CM12_29 node13_3 node13_8 -3.878491e-15
CM12_30 node13_3 node13_9 -4.144789e-15
CM12_31 node13_4 node13_5 -3.011387e-13
CM12_32 node13_4 node13_6 -2.590566e-14
CM12_33 node13_4 node13_7 -1.142857e-14
CM12_34 node13_4 node13_8 -6.642276e-15
CM12_35 node13_4 node13_9 -6.914501e-15
CM12_36 node13_5 node13_6 -3.012291e-13
CM12_37 node13_5 node13_7 -2.628136e-14
CM12_38 node13_5 node13_8 -1.220907e-14
CM12_39 node13_5 node13_9 -1.177964e-14
CM12_40 node13_6 node13_7 -3.018016e-13
CM12_41 node13_6 node13_8 -2.762580e-14
CM12_42 node13_6 node13_9 -2.099353e-14
CM12_43 node13_7 node13_8 -3.042640e-13
CM12_44 node13_7 node13_9 -4.332676e-14
CM12_45 node13_8 node13_9 -3.372029e-13
R13_1 node13_0 node13_0_mid 6.559697e-02
L13_1 node13_0_mid node14_0 1.324593e-01
R13_2 node13_1 node13_1_mid 6.559697e-02
L13_2 node13_1_mid node14_1 1.324593e-01
R13_3 node13_2 node13_2_mid 6.559697e-02
L13_3 node13_2_mid node14_2 1.324592e-01
R13_4 node13_3 node13_3_mid 6.559697e-02
L13_4 node13_3_mid node14_3 1.324592e-01
R13_5 node13_4 node13_4_mid 6.559697e-02
L13_5 node13_4_mid node14_4 1.324592e-01
R13_6 node13_5 node13_5_mid 6.559697e-02
L13_6 node13_5_mid node14_5 1.324591e-01
R13_7 node13_6 node13_6_mid 6.559697e-02
L13_7 node13_6_mid node14_6 1.324591e-01
R13_8 node13_7 node13_7_mid 6.559697e-02
L13_8 node13_7_mid node14_7 1.324591e-01
R13_9 node13_8 node13_8_mid 6.559697e-02
L13_9 node13_8_mid node14_8 1.324591e-01
R13_10 node13_9 node13_9_mid 6.559697e-02
L13_10 node13_9_mid node14_9 1.324591e-01
K13_1 L13_1 L13_2 1.000000e+00
K13_2 L13_1 L13_3 1.000000e+00
K13_3 L13_1 L13_4 1.000000e+00
K13_4 L13_1 L13_5 1.000000e+00
K13_5 L13_1 L13_6 9.999999e-01
K13_6 L13_1 L13_7 1.000000e+00
K13_7 L13_1 L13_8 9.999999e-01
K13_8 L13_1 L13_9 9.999999e-01
K13_9 L13_1 L13_10 9.999999e-01
K13_10 L13_2 L13_3 1.000000e+00
K13_11 L13_2 L13_4 1.000000e+00
K13_12 L13_2 L13_5 1.000000e+00
K13_13 L13_2 L13_6 9.999999e-01
K13_14 L13_2 L13_7 1.000000e+00
K13_15 L13_2 L13_8 9.999999e-01
K13_16 L13_2 L13_9 9.999999e-01
K13_17 L13_2 L13_10 9.999999e-01
K13_18 L13_3 L13_4 1.000000e+00
K13_19 L13_3 L13_5 1.000000e+00
K13_20 L13_3 L13_6 9.999999e-01
K13_21 L13_3 L13_7 9.999999e-01
K13_22 L13_3 L13_8 9.999999e-01
K13_23 L13_3 L13_9 9.999999e-01
K13_24 L13_3 L13_10 9.999998e-01
K13_25 L13_4 L13_5 1.000000e+00
K13_26 L13_4 L13_6 9.999999e-01
K13_27 L13_4 L13_7 1.000000e+00
K13_28 L13_4 L13_8 9.999999e-01
K13_29 L13_4 L13_9 9.999999e-01
K13_30 L13_4 L13_10 9.999999e-01
K13_31 L13_5 L13_6 9.999999e-01
K13_32 L13_5 L13_7 1.000000e+00
K13_33 L13_5 L13_8 9.999999e-01
K13_34 L13_5 L13_9 9.999999e-01
K13_35 L13_5 L13_10 9.999999e-01
K13_36 L13_6 L13_7 9.999999e-01
K13_37 L13_6 L13_8 1.000000e+00
K13_38 L13_6 L13_9 1.000000e+00
K13_39 L13_6 L13_10 9.999999e-01
K13_40 L13_7 L13_8 9.999999e-01
K13_41 L13_7 L13_9 9.999999e-01
K13_42 L13_7 L13_10 9.999999e-01
K13_43 L13_8 L13_9 1.000000e+00
K13_44 L13_8 L13_10 1.000000e+00
K13_45 L13_9 L13_10 1.000000e+00
C13_1 node14_0 0 4.303416e-13
G13_1 node14_0 0 node14_0 0 2.703916e-06
C13_2 node14_1 0 6.975560e-13
G13_2 node14_1 0 node14_1 0 4.382874e-06
C13_3 node14_2 0 7.023171e-13
G13_3 node14_2 0 node14_2 0 4.412789e-06
C13_4 node14_3 0 7.031524e-13
G13_4 node14_3 0 node14_3 0 4.418037e-06
C13_5 node14_4 0 7.034466e-13
G13_5 node14_4 0 node14_4 0 4.419885e-06
C13_6 node14_5 0 7.035676e-13
G13_6 node14_5 0 node14_5 0 4.420645e-06
C13_7 node14_6 0 7.030741e-13
G13_7 node14_6 0 node14_6 0 4.417545e-06
C13_8 node14_7 0 7.018853e-13
G13_8 node14_7 0 node14_7 0 4.410075e-06
C13_9 node14_8 0 6.973380e-13
G13_9 node14_8 0 node14_8 0 4.381504e-06
C13_10 node14_9 0 4.303249e-13
G13_10 node14_9 0 node14_9 0 2.703811e-06
CM13_1 node14_0 node14_1 -3.372270e-13
CM13_2 node14_0 node14_2 -4.333637e-14
CM13_3 node14_0 node14_3 -2.097687e-14
CM13_4 node14_0 node14_4 -1.177420e-14
CM13_5 node14_0 node14_5 -6.918544e-15
CM13_6 node14_0 node14_6 -4.146150e-15
CM13_7 node14_0 node14_7 -2.537949e-15
CM13_8 node14_0 node14_8 -1.643541e-15
CM13_9 node14_0 node14_9 -1.780983e-15
CM13_10 node14_1 node14_2 -3.044883e-13
CM13_11 node14_1 node14_3 -2.759806e-14
CM13_12 node14_1 node14_4 -1.220281e-14
CM13_13 node14_1 node14_5 -6.645893e-15
CM13_14 node14_1 node14_6 -3.879486e-15
CM13_15 node14_1 node14_7 -2.352696e-15
CM13_16 node14_1 node14_8 -1.518489e-15
CM13_17 node14_1 node14_9 -1.643380e-15
CM13_18 node14_2 node14_3 -3.019823e-13
CM13_19 node14_2 node14_4 -2.628447e-14
CM13_20 node14_2 node14_5 -1.143815e-14
CM13_21 node14_2 node14_6 -6.217217e-15
CM13_22 node14_2 node14_7 -3.678469e-15
CM13_23 node14_2 node14_8 -2.353400e-15
CM13_24 node14_2 node14_9 -2.538483e-15
CM13_25 node14_3 node14_4 -3.011554e-13
CM13_26 node14_3 node14_5 -2.592703e-14
CM13_27 node14_3 node14_6 -1.127554e-14
CM13_28 node14_3 node14_7 -6.213871e-15
CM13_29 node14_3 node14_8 -3.878491e-15
CM13_30 node14_3 node14_9 -4.144789e-15
CM13_31 node14_4 node14_5 -3.011387e-13
CM13_32 node14_4 node14_6 -2.590566e-14
CM13_33 node14_4 node14_7 -1.142857e-14
CM13_34 node14_4 node14_8 -6.642276e-15
CM13_35 node14_4 node14_9 -6.914501e-15
CM13_36 node14_5 node14_6 -3.012291e-13
CM13_37 node14_5 node14_7 -2.628136e-14
CM13_38 node14_5 node14_8 -1.220907e-14
CM13_39 node14_5 node14_9 -1.177964e-14
CM13_40 node14_6 node14_7 -3.018016e-13
CM13_41 node14_6 node14_8 -2.762580e-14
CM13_42 node14_6 node14_9 -2.099353e-14
CM13_43 node14_7 node14_8 -3.042640e-13
CM13_44 node14_7 node14_9 -4.332676e-14
CM13_45 node14_8 node14_9 -3.372029e-13
R_in1 in1 node0_0 1e-6
R_out1 node14_0 out1 1e-6
R_in2 in2 node0_1 1e-6
R_out2 node14_1 out2 1e-6
R_in3 in3 node0_2 1e-6
R_out3 node14_2 out3 1e-6
R_in4 in4 node0_3 1e-6
R_out4 node14_3 out4 1e-6
R_in5 in5 node0_4 1e-6
R_out5 node14_4 out5 1e-6
R_in6 in6 node0_5 1e-6
R_out6 node14_5 out6 1e-6
R_in7 in7 node0_6 1e-6
R_out7 node14_6 out7 1e-6
R_in8 in8 node0_7 1e-6
R_out8 node14_7 out8 1e-6
R_in9 in9 node0_8 1e-6
R_out9 node14_8 out9 1e-6
R_in10 in10 node0_9 1e-6
R_out10 node14_9 out10 1e-6
.ENDS TRANSMISSION_LINE
