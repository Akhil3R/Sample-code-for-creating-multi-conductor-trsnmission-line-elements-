* 10-wire PI Transmission Line Subcircuit Model

.SUBCKT TRANSMISSION_LINE in1 out1 in2 out2 in3 out3 in4 out4 in5 out5 in6 out6 in7 out7 in8 out8 in9 out9 in10 out10 
R0_1 node0_0 node0_0_mid 6.887682e-02
L0_1 node0_0_mid node1_0 1.390822e-01
R0_2 node0_1 node0_1_mid 6.887682e-02
L0_2 node0_1_mid node1_1 1.390822e-01
R0_3 node0_2 node0_2_mid 6.887682e-02
L0_3 node0_2_mid node1_2 1.390822e-01
R0_4 node0_3 node0_3_mid 6.887682e-02
L0_4 node0_3_mid node1_3 1.390821e-01
R0_5 node0_4 node0_4_mid 6.887682e-02
L0_5 node0_4_mid node1_4 1.390821e-01
R0_6 node0_5 node0_5_mid 6.887682e-02
L0_6 node0_5_mid node1_5 1.390821e-01
R0_7 node0_6 node0_6_mid 6.887682e-02
L0_7 node0_6_mid node1_6 1.390820e-01
R0_8 node0_7 node0_7_mid 6.887682e-02
L0_8 node0_7_mid node1_7 1.390820e-01
R0_9 node0_8 node0_8_mid 6.887682e-02
L0_9 node0_8_mid node1_8 1.390820e-01
R0_10 node0_9 node0_9_mid 6.887682e-02
L0_10 node0_9_mid node1_9 1.390821e-01
K0_1 L0_1 L0_2 1.000000e+00
K0_2 L0_1 L0_3 1.000000e+00
K0_3 L0_1 L0_4 1.000000e+00
K0_4 L0_1 L0_5 1.000000e+00
K0_5 L0_1 L0_6 9.999999e-01
K0_6 L0_1 L0_7 1.000000e+00
K0_7 L0_1 L0_8 9.999999e-01
K0_8 L0_1 L0_9 9.999999e-01
K0_9 L0_1 L0_10 9.999999e-01
K0_10 L0_2 L0_3 1.000000e+00
K0_11 L0_2 L0_4 1.000000e+00
K0_12 L0_2 L0_5 1.000000e+00
K0_13 L0_2 L0_6 9.999999e-01
K0_14 L0_2 L0_7 1.000000e+00
K0_15 L0_2 L0_8 9.999999e-01
K0_16 L0_2 L0_9 9.999999e-01
K0_17 L0_2 L0_10 9.999999e-01
K0_18 L0_3 L0_4 1.000000e+00
K0_19 L0_3 L0_5 1.000000e+00
K0_20 L0_3 L0_6 9.999999e-01
K0_21 L0_3 L0_7 9.999999e-01
K0_22 L0_3 L0_8 9.999999e-01
K0_23 L0_3 L0_9 9.999999e-01
K0_24 L0_3 L0_10 9.999998e-01
K0_25 L0_4 L0_5 1.000000e+00
K0_26 L0_4 L0_6 9.999999e-01
K0_27 L0_4 L0_7 1.000000e+00
K0_28 L0_4 L0_8 9.999999e-01
K0_29 L0_4 L0_9 9.999999e-01
K0_30 L0_4 L0_10 9.999999e-01
K0_31 L0_5 L0_6 9.999999e-01
K0_32 L0_5 L0_7 1.000000e+00
K0_33 L0_5 L0_8 9.999999e-01
K0_34 L0_5 L0_9 9.999999e-01
K0_35 L0_5 L0_10 9.999999e-01
K0_36 L0_6 L0_7 9.999999e-01
K0_37 L0_6 L0_8 1.000000e+00
K0_38 L0_6 L0_9 1.000000e+00
K0_39 L0_6 L0_10 9.999999e-01
K0_40 L0_7 L0_8 9.999999e-01
K0_41 L0_7 L0_9 9.999999e-01
K0_42 L0_7 L0_10 9.999999e-01
K0_43 L0_8 L0_9 1.000000e+00
K0_44 L0_8 L0_10 1.000000e+00
K0_45 L0_9 L0_10 1.000000e+00
C0_1 node1_0 0 4.518586e-13
G0_1 node1_0 0 node1_0 0 2.839112e-06
C0_2 node1_1 0 7.324338e-13
G0_2 node1_1 0 node1_1 0 4.602017e-06
C0_3 node1_2 0 7.374330e-13
G0_3 node1_2 0 node1_2 0 4.633428e-06
C0_4 node1_3 0 7.383100e-13
G0_4 node1_3 0 node1_3 0 4.638939e-06
C0_5 node1_4 0 7.386189e-13
G0_5 node1_4 0 node1_4 0 4.640879e-06
C0_6 node1_5 0 7.387459e-13
G0_6 node1_5 0 node1_5 0 4.641678e-06
C0_7 node1_6 0 7.382278e-13
G0_7 node1_6 0 node1_6 0 4.638422e-06
C0_8 node1_7 0 7.369795e-13
G0_8 node1_7 0 node1_7 0 4.630579e-06
C0_9 node1_8 0 7.322049e-13
G0_9 node1_8 0 node1_8 0 4.600579e-06
C0_10 node1_9 0 4.518411e-13
G0_10 node1_9 0 node1_9 0 2.839001e-06
CM0_1 node1_0 node1_1 -3.540883e-13
CM0_2 node1_0 node1_2 -4.550319e-14
CM0_3 node1_0 node1_3 -2.202572e-14
CM0_4 node1_0 node1_4 -1.236291e-14
CM0_5 node1_0 node1_5 -7.264472e-15
CM0_6 node1_0 node1_6 -4.353458e-15
CM0_7 node1_0 node1_7 -2.664846e-15
CM0_8 node1_0 node1_8 -1.725718e-15
CM0_9 node1_0 node1_9 -1.870032e-15
CM0_10 node1_1 node1_2 -3.197127e-13
CM0_11 node1_1 node1_3 -2.897796e-14
CM0_12 node1_1 node1_4 -1.281295e-14
CM0_13 node1_1 node1_5 -6.978188e-15
CM0_14 node1_1 node1_6 -4.073460e-15
CM0_15 node1_1 node1_7 -2.470330e-15
CM0_16 node1_1 node1_8 -1.594413e-15
CM0_17 node1_1 node1_9 -1.725549e-15
CM0_18 node1_2 node1_3 -3.170814e-13
CM0_19 node1_2 node1_4 -2.759870e-14
CM0_20 node1_2 node1_5 -1.201006e-14
CM0_21 node1_2 node1_6 -6.528078e-15
CM0_22 node1_2 node1_7 -3.862392e-15
CM0_23 node1_2 node1_8 -2.471070e-15
CM0_24 node1_2 node1_9 -2.665407e-15
CM0_25 node1_3 node1_4 -3.162132e-13
CM0_26 node1_3 node1_5 -2.722338e-14
CM0_27 node1_3 node1_6 -1.183931e-14
CM0_28 node1_3 node1_7 -6.524565e-15
CM0_29 node1_3 node1_8 -4.072416e-15
CM0_30 node1_3 node1_9 -4.352028e-15
CM0_31 node1_4 node1_5 -3.161957e-13
CM0_32 node1_4 node1_6 -2.720094e-14
CM0_33 node1_4 node1_7 -1.200000e-14
CM0_34 node1_4 node1_8 -6.974389e-15
CM0_35 node1_4 node1_9 -7.260226e-15
CM0_36 node1_5 node1_6 -3.162906e-13
CM0_37 node1_5 node1_7 -2.759542e-14
CM0_38 node1_5 node1_8 -1.281953e-14
CM0_39 node1_5 node1_9 -1.236862e-14
CM0_40 node1_6 node1_7 -3.168916e-13
CM0_41 node1_6 node1_8 -2.900709e-14
CM0_42 node1_6 node1_9 -2.204321e-14
CM0_43 node1_7 node1_8 -3.194772e-13
CM0_44 node1_7 node1_9 -4.549309e-14
CM0_45 node1_8 node1_9 -3.540630e-13
R_in1 in1 node0_0 1e-6
R_out1 node1_0 out1 1e-6
R_in2 in2 node0_1 1e-6
R_out2 node1_1 out2 1e-6
R_in3 in3 node0_2 1e-6
R_out3 node1_2 out3 1e-6
R_in4 in4 node0_3 1e-6
R_out4 node1_3 out4 1e-6
R_in5 in5 node0_4 1e-6
R_out5 node1_4 out5 1e-6
R_in6 in6 node0_5 1e-6
R_out6 node1_5 out6 1e-6
R_in7 in7 node0_6 1e-6
R_out7 node1_6 out7 1e-6
R_in8 in8 node0_7 1e-6
R_out8 node1_7 out8 1e-6
R_in9 in9 node0_8 1e-6
R_out9 node1_8 out9 1e-6
R_in10 in10 node0_9 1e-6
R_out10 node1_9 out10 1e-6
.ENDS TRANSMISSION_LINE
